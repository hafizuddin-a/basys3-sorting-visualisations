`timescale 1ns / 1ps

module top_module (
    input btnC,
    input btnU,
    input btnD, 
    input btnL, 
    input btnR,
    input [0:15] sw,
    output reg [15:0] led = 0,
    
    input clk,
    output [7:0] Jx,
    output [7:0] JXADC,
    output reg [0:3] an = 4'b1111,
    output reg [0:6] seg = 7'b1111111
);

    wire frame_begin, sending_pixels, sample_pixel;
    wire frame_begin2, sending_pixels2, sample_pixel2;    
    wire [12:0] pixel_index;
    wire [12:0] pixel_index2;
    reg [15:0] oled_data;
    reg [15:0] oled_data2;
    wire clk_6p25m;
    
    // 7 seg display 
    reg [16:0] seven_seg_counter = 0;
    reg [1:0] anode_index = 0;
    reg [3:0] sorting_algorithm = 0; // 0001 = bubble; 0010 = selection; 0100 = insertion; 1000 = cocktail; 0011 = dOnE
    
    clk6p25m clock_display(clk, clk_6p25m);
    
    Oled_Display unit_oled (
        .clk(clk_6p25m), 
        .reset(0), 
        .frame_begin(frame_begin), 
        .sending_pixels(sending_pixels),
        .sample_pixel(sample_pixel), 
        .pixel_index(pixel_index), 
        .pixel_data(oled_data), 
        .cs(Jx[0]), 
        .sdin(Jx[1]), 
        .sclk(Jx[3]), 
        .d_cn(Jx[4]), 
        .resn(Jx[5]), 
        .vccen(Jx[6]), 
        .pmoden(Jx[7])
    );
    
    Oled_Display unit_oled2 (
        .clk(clk_6p25m), 
        .reset(0), 
        .frame_begin(frame_begin2), 
        .sending_pixels(sending_pixels2),
        .sample_pixel(sample_pixel2), 
        .pixel_index(pixel_index2), 
        .pixel_data(oled_data2), 
        .cs(JXADC[0]), 
        .sdin(JXADC[1]), 
        .sclk(JXADC[3]), 
        .d_cn(JXADC[4]), 
        .resn(JXADC[5]), 
        .vccen(JXADC[6]), 
        .pmoden(JXADC[7])
    );
     
    // Parameters for bar display
    localparam BAR_WIDTH = 8;
    localparam BAR_SPACING = 2;
    localparam BAR_COLOR = 16'h07E0; // Green color
    localparam BACKGROUND_COLOR = 16'h0000; // Black background
    localparam SORT_DELAY = 100_000_000; // Delay between sort steps (adjust as needed)
    
    reg [6:0] key;
    reg [6:0] bar_heights [4:0];
    reg [6:0] counter;
    reg [31:0] delay_counter; // Counter for sorting delay
    reg sorting = 0; // Flag to indicate sorting is in progress
    reg [4:0] is_bar_sorted = 5'b00000; // If true, green; yellow otherwise
    reg sorted; // Flag to indicate sorting is complete
    integer i, j, k, min_index;
    reg dir; // Flag for direction of sorting
    reg random_bars_generated;
    reg [3:0] curr_digit_manual; // Digit to manually input from 1 - 9
    reg [2:0] curr_index_manual = 3'b000; // Digit index for manual input
    wire btnC_debouncer;
    reg is_finished_manual_input = 0;
    debouncer centre_debouncer(clk, btnC, btnC_debouncer);
    reg is_begin_manual_input = 0;
    reg [23:0] looping_counter = 0;
    reg [4:0] looping_leds = 1;
    reg [3:0] looping_7_seg = 0;
    integer movement = 0;
    reg swap;
    integer swap_from = 10;
    integer swap_to = 10;
    integer selection_sort_from;
    integer selection_sort_to;
    
    // 2nd OLED
    reg [31:0] menucounter = 0; // Counter to keep track of clock cycles
    reg [2:0] menuframe = 0; // Register to store the current frame
    reg [31:0] celebcounter = 0;
    reg [5:0] celebframe = 1;

    always @ (posedge clk) begin 

        sorting_algorithm = btnU ? 4'b0001 : 
                            btnD ? 4'b0010 : 
                            btnR ? 4'b0100 : 
                            btnL ? 4'b1000 : sorting_algorithm;
                            
        // Frame count for main menu
        if (sorting_algorithm == 0 || sorting_algorithm == 4'b0011) begin
            menucounter <= menucounter + 1; // Increment counter on every clock cycle
            celebcounter <= celebcounter + 1;
    
            
            if (menucounter == 100000000) begin
                menucounter <= 0; // Reset counter
                menuframe <= (menuframe == 6) ? 0 : menuframe + 1; // Increment frame or reset to 0 if at frame 7 
            end
            
            if (celebcounter == 10000000) begin
                celebcounter <= 0; // Reset counter
                celebframe <= (celebframe == 12) ? 1 : celebframe + 1;
            end
	end
        
        seven_seg_counter <= seven_seg_counter + 1;
        looping_counter <= looping_counter + 1;
        if (seven_seg_counter == 100_000) begin 
            seven_seg_counter <= 0;
            anode_index <= anode_index + 1;
        end
        
        if (looping_counter == 10_000_000) begin
            looping_counter <= 0;
        end
        
        if (sw[15]) begin // Reset
            bar_heights[0] = 0;
            bar_heights[1] = 0;
            bar_heights[2] = 0;
            bar_heights[3] = 0;
            bar_heights[4] = 0;
            random_bars_generated <= 0;
            is_begin_manual_input <= 0;
            sorting <= 0;
            is_finished_manual_input <= 0;
            sorted <= 0;
            curr_index_manual <= 0;
            led <= 0;
            seg <= 7'b1111111;
            an <= 4'b1111;
            sorting_algorithm <= 4'b0000;
        end
        
        if (sorting_algorithm == 4'b0001) begin // Bubble sort
            case (anode_index) 
                2'b00: begin 
                    an = 4'b0111;
                    seg = 7'b1110001;
                end
                2'b01: begin 
                    an = 4'b1011;
                    seg = 7'b1100000;
                end
                2'b10: begin 
                    an = 4'b1101;
                    seg = 7'b1000001;
                end
                2'b11: begin 
                    an = 4'b1110;
                    seg = 7'b1100000;
                end
            endcase
            if (!is_begin_manual_input && btnC_debouncer && !sorting) begin 
                is_begin_manual_input = 1;
            end else if (!sw[0] && !is_finished_manual_input && is_begin_manual_input) begin // Manual input mode 
                sorting <= 0;
                delay_counter <= 0;
                j <= 0;
                random_bars_generated <= 0; // Reset the flag
                sorted <= 0; // Reset the sorted flag
                if (!btnC && curr_index_manual < 5) begin 
                    curr_digit_manual = sw[9] ? 9 : sw[8] ? 8 : sw[7] ? 7 : sw[6] ? 6 : sw[5] ? 5 :
                                        sw[4] ? 4 : sw[3] ? 3 : sw[2] ? 2 : sw[1] ? 1 : 1;
                    bar_heights[curr_index_manual] <= curr_digit_manual * 7;
                    if (curr_index_manual < 5 ) 
                        led[curr_index_manual] <= 1;
                end else begin
                    if (curr_index_manual == 5) 
                        curr_index_manual <= 0;
                    if (btnC_debouncer) begin 
                        led[curr_index_manual] <= 1;
                        curr_index_manual <= curr_index_manual + 1;
                        if (curr_index_manual == 5) 
                            is_finished_manual_input <= 1;
                            is_begin_manual_input <= 0;
                    end
                end
            end else if (sw[0] && !btnU && !random_bars_generated) begin // Random input mode
                counter <= counter + 1; // Increment counter
                is_finished_manual_input = 0;
                for (i = 0; i < 5; i = i + 1) begin
                    bar_heights[i] <= (counter * 37 + i * 17) % 63 + 1; // Generate more random heights
                end
                sorting <= 0; // Ensure sorting is not started yet
                delay_counter <= 0;
                j <= 0;
                random_bars_generated <= 1; // Set the flag
                sorted <= 0; // Reset the sorted flag
                
            end else if (btnU && !sorting && !sorted && (is_finished_manual_input || random_bars_generated)) begin
                sorting <= 1; // Start sorting
                i <= 0; // Initialize indices for bubble sort
                j <= 0;
            end else if (sorting) begin // Bubble sort
                led[5:0] <= looping_leds; // Loading led
                if (looping_counter == 0) begin
                    looping_leds <= {looping_leds[3:0], looping_leds[4]};
                    looping_7_seg <= (looping_7_seg == 11) ? 0 : looping_7_seg + 1;
                end
                case (looping_7_seg) // Loading 7-seg
                    0: begin
                        an = 4'b0111;
                        seg = 7'b0111111;
                    end
                    1: begin
                        an = 4'b0111;
                        seg = 7'b1011111;
                    end
                    2: begin
                        an = 4'b0111;
                        seg = 7'b1101111;
                    end
                    3: begin
                        an = 4'b0111;
                        seg = 7'b1110111;
                    end
                    4: begin
                        an = 4'b1011;
                        seg = 7'b1110111;
                    end
                    5: begin
                        an = 4'b1101;
                        seg = 7'b1110111;
                    end
                    6: begin
                        an = 4'b1110;
                        seg = 7'b1110111;
                    end
                    7: begin
                        an = 4'b1110;
                        seg = 7'b1111011;
                    end
                    8: begin
                        an = 4'b1110;
                        seg = 7'b1111101;
                    end
                    9: begin
                        an = 4'b1110;
                        seg = 7'b0111111;
                    end
                    10: begin
                        an = 4'b1101;
                        seg = 7'b0111111;
                    end
                    11: begin
                        an = 4'b1011;
                        seg = 7'b0111111;
                    end
                endcase
                if (delay_counter < SORT_DELAY) begin
                    delay_counter <= delay_counter + 1; // Increment delay counter
                end else begin
                    delay_counter <= 0; // Reset delay counter
                    if (j < 4 - i) begin
                        if (bar_heights[j] > bar_heights[j + 1]) begin
                            // Swap adjacent bars if they are in the wrong order
                            {bar_heights[j], bar_heights[j + 1]} <= {bar_heights[j + 1], bar_heights[j]};
                            swap_from <= j;
                            swap_to <= j + 1;
                            swap <= 1;
                        end else begin
                            swap_from <= 10;
                            swap_to <= 10; 
                            swap <= 0;
                        end
                        j <= j + 1; // Move to the next pair
                    end else begin
                        swap_from <= 10;
                        swap_to <= 10; 
                        swap <= 0;
                        if (i < 3) begin
                            i <= i + 1; // Move to the next pass of the bubble sort
                            j <= 0; // Reset the inner loop counter
                        end else begin
                            sorting <= 0; // Sorting is complete
                            sorted <= 1; // Set the sorted flag
                            is_begin_manual_input <= 0;
                            sorting_algorithm <= 4'b0011; // Display dOnE
                        end
                    end
                end
            end
        end
        
        else if (sorting_algorithm == 4'b0010) begin // Selection sort
            case (anode_index) 
                2'b00: begin
                    an = 4'b0111;
                    seg = 7'b0110001;
                end
                2'b01: begin
                    an = 4'b1011;
                    seg = 7'b1110001;
                end
                2'b10: begin
                    an = 4'b1101;
                    seg = 7'b0110000;
                end
                2'b11: begin
                    an = 4'b1110;
                    seg = 7'b0100100;
                end
            endcase
            if (!is_begin_manual_input && btnC_debouncer && !sorting) begin 
                is_begin_manual_input = 1;
            end else if (!sw[0] && !is_finished_manual_input) begin // Manual input mode 
                sorting <= 0;
                delay_counter <= 0;
                j <= 0;
                random_bars_generated <= 0; // Reset the flag
                sorted <= 0; // Reset the sorted flag
                if (!btnC && curr_index_manual < 5) begin 
                    curr_digit_manual = sw[9] ? 9 : sw[8] ? 8 : sw[7] ? 7 : sw[6] ? 6 : sw[5] ? 5 :
                                        sw[4] ? 4 : sw[3] ? 3 : sw[2] ? 2 : sw[1] ? 1 : 1;
                    bar_heights[curr_index_manual] <= curr_digit_manual * 7;
                    led[curr_index_manual] <= 1;
                end else if (btnC_debouncer) begin
                    led[curr_index_manual] <= 1;
                    curr_index_manual <= curr_index_manual + 1;
                    if (curr_index_manual == 5) 
                        is_finished_manual_input <= 1;
                end
            end else if (sw[0] && !btnD && !random_bars_generated) begin // Random input mode
                counter <= counter + 1; // Increment counter
                is_finished_manual_input = 0;
                for (i = 0; i < 5; i = i + 1) begin
                    bar_heights[i] <= (counter * 37 + i * 17) % 63 + 1; // Generate more random heights
                end
                sorting <= 0; // Ensure sorting is not started yet
                delay_counter <= 0;
                j <= 0;
                random_bars_generated <= 1; // Set the flag
                sorted <= 0; // Reset the sorted flag
            end else if (btnD && !sorting && !sorted && (is_finished_manual_input || random_bars_generated)) begin
                sorting <= 1; // Start sorting
                i <= 0; // Initialize indices for bubble sort
                j <= 0;
                min_index <= i; // Set min_index to i for the first pass
            end else if (sorting && !sorted) begin // Selection sort
                led[5:0] <= looping_leds; // Loading led
                if (looping_counter == 0) begin
                    looping_leds <= {looping_leds[3:0], looping_leds[4]};
                    looping_7_seg <= (looping_7_seg == 11) ? 0 : looping_7_seg + 1;
                end
                case (looping_7_seg) // Loading 7-seg
                    0: begin
                        an = 4'b0111;
                        seg = 7'b0111111;
                    end
                    1: begin
                        an = 4'b0111;
                        seg = 7'b1011111;
                    end
                    2: begin
                        an = 4'b0111;
                        seg = 7'b1101111;
                    end
                    3: begin
                        an = 4'b0111;
                        seg = 7'b1110111;
                    end
                    4: begin
                        an = 4'b1011;
                        seg = 7'b1110111;
                    end
                    5: begin
                        an = 4'b1101;
                        seg = 7'b1110111;
                    end
                    6: begin
                        an = 4'b1110;
                        seg = 7'b1110111;
                    end
                    7: begin
                        an = 4'b1110;
                        seg = 7'b1111011;
                    end
                    8: begin
                        an = 4'b1110;
                        seg = 7'b1111101;
                    end
                    9: begin
                        an = 4'b1110;
                        seg = 7'b0111111;
                    end
                    10: begin
                        an = 4'b1101;
                        seg = 7'b0111111;
                    end
                    11: begin
                        an = 4'b1011;
                        seg = 7'b0111111;
                    end
                endcase  
                if (delay_counter < SORT_DELAY) begin
                    delay_counter <= delay_counter + 1; // Increment delay counter
                end else begin
                    delay_counter <= 0; // Reset delay counter
                    if (i < 5) begin // Change condition to iterate for all 5 passes
                        if (j < 5) begin
                            if (j > i) begin
                                if (bar_heights[j] < bar_heights[min_index]) begin
                                    min_index <= j; // Update the index of the minimum value
                                end
                            end
                            j <= j + 1; // Move to the next index
                            swap_from <= 10;
                            swap_to <= 10;
                            swap <= 0;
                        end else begin
                            // Swap the values at i and min_index
                            if (min_index != i) begin
                                {bar_heights[i], bar_heights[min_index]} <= {bar_heights[min_index], bar_heights[i]}; 
                            end
                            i <= i + 1; // Move to the next pass of the selection sort
                            j <= i + 1; // Reset inner loop counter
                            min_index <= i + 1; // Reset min_index
                        end
                    end else begin
                        sorting <= 0; // Sorting is complete
                        sorted <= 1; // Set sorted flag
                        is_finished_manual_input <= 0;
                        sorting_algorithm <= 4'b0011; // Display dOnE
                        i <= 0;
                        j <= 0;
                    end
                end
            end
        end
        
        else if (sorting_algorithm == 4'b0100) begin // Insertion sort
            case (anode_index) 
                2'b00: begin
                    an = 4'b0111;
                    seg = 7'b1111010;
                end
                2'b01: begin
                    an = 4'b1011;
                    seg = 7'b0100100;
                end
                2'b10: begin
                    an = 4'b1101;
                    seg = 7'b1101010;
                end
                2'b11: begin
                    an = 4'b1110;
                    seg = 7'b1001111;
                end
            endcase
            if (!is_begin_manual_input && btnC_debouncer && !sorting) begin 
                is_begin_manual_input = 1;
            end else if (!sw[0] && !is_finished_manual_input) begin // Manual input mode 
                sorting <= 0;
                delay_counter <= 0;
                j <= 0;
                random_bars_generated <= 0; // Reset the flag
                sorted <= 0; // Reset the sorted flag
                is_bar_sorted <= 0;
                if (!btnC && curr_index_manual < 5) begin 
                    curr_digit_manual = sw[9] ? 9 : sw[8] ? 8 : sw[7] ? 7 : sw[6] ? 6 : sw[5] ? 5 :
                                        sw[4] ? 4 : sw[3] ? 3 : sw[2] ? 2 : sw[1] ? 1 : 1;
                    bar_heights[curr_index_manual] <= curr_digit_manual * 7;
                    led[curr_index_manual] <= 1;
                end else if (btnC_debouncer) begin
                    led[curr_index_manual] <= 1;
                    curr_index_manual <= curr_index_manual + 1;
                    if (curr_index_manual == 5) 
                        is_finished_manual_input <= 1;
                end
            end else if (sw[0] && !btnR && !random_bars_generated) begin // Random input mode
                counter <= counter + 1; // Increment counter
                is_finished_manual_input = 0;
                for (i = 0; i < 5; i = i + 1) begin
                    bar_heights[i] <= (counter * 37 + i * 17) % 63 + 1; // Generate more random heights
                end
                sorting <= 0; // Ensure sorting is not started yet
                delay_counter <= 0;
                j <= 0;
                random_bars_generated <= 1; // Set the flag
                sorted <= 0; // Reset the sorted flag
            end else if (btnR && !sorting && !sorted && (is_finished_manual_input || random_bars_generated)) begin
                sorting <= 1; // Start sorting
                i <= 1; // Initialize indices for bubble sort
                j <= 1;
                is_bar_sorted <= 5'b10000;
            end else if (sorting) begin // Insertion sort
                led[5:0] <= looping_leds; // Loading led
                if (looping_counter == 0) begin
                    looping_leds <= {looping_leds[3:0], looping_leds[4]};
                    looping_7_seg <= (looping_7_seg == 11) ? 0 : looping_7_seg + 1;
                end
                case (looping_7_seg) // Loading 7-seg
                    0: begin
                        an = 4'b0111;
                        seg = 7'b0111111;
                    end
                    1: begin
                        an = 4'b0111;
                        seg = 7'b1011111;
                    end
                    2: begin
                        an = 4'b0111;
                        seg = 7'b1101111;
                    end
                    3: begin
                        an = 4'b0111;
                        seg = 7'b1110111;
                    end
                    4: begin
                        an = 4'b1011;
                        seg = 7'b1110111;
                    end
                    5: begin
                        an = 4'b1101;
                        seg = 7'b1110111;
                    end
                    6: begin
                        an = 4'b1110;
                        seg = 7'b1110111;
                    end
                    7: begin
                        an = 4'b1110;
                        seg = 7'b1111011;
                    end
                    8: begin
                        an = 4'b1110;
                        seg = 7'b1111101;
                    end
                    9: begin
                        an = 4'b1110;
                        seg = 7'b0111111;
                    end
                    10: begin
                        an = 4'b1101;
                        seg = 7'b0111111;
                    end
                    11: begin
                        an = 4'b1011;
                        seg = 7'b0111111;
                    end
                endcase  
                if (delay_counter < SORT_DELAY) begin
                    delay_counter <= delay_counter + 1; // Increment delay counter
                end else begin
                    delay_counter <= 0; // Reset delay counter
                    if (i < 4) begin
                        if (j >= 0 && bar_heights[j + 1] < bar_heights[j]) begin //CHANGE HERE?
                            {bar_heights[j + 1], bar_heights[j]} <= {bar_heights[j], bar_heights[j + 1]};
                            swap_from <= j;
                            swap_to <= j + 1; 
                            swap <= 1;
                            j <= j - 1;
                        end else begin
                            swap_from <= 10;
                            swap_to <= 10; 
                            swap <= 0;
                            case (i)
                            0: is_bar_sorted <= is_bar_sorted + 5'b01000;
                            1: is_bar_sorted <= is_bar_sorted + 5'b00100;
                            2: is_bar_sorted <= is_bar_sorted + 5'b00010;
                            3: is_bar_sorted <= is_bar_sorted + 5'b00001;
                            endcase
                            i = i + 1;
                            j = i;
                        end
                    end else begin 
                        sorted <= 1;
                        sorting <= 0;
                        is_finished_manual_input <= 0;
                        sorting_algorithm <= 4'b0011; // Display dOnE
                    end
                end
            end
        end
        
        else if (sorting_algorithm == 4'b1000) begin // Cocktail sort
            case (anode_index) 
                2'b00: begin
                    an = 4'b0111;
                    seg = 7'b1010000;
                end
                2'b01: begin
                    an = 4'b1011;
                    seg = 7'b0110001;
                end
                2'b10: begin
                    an = 4'b1101;
                    seg = 7'b0000001;
                end
                2'b11: begin
                    an = 4'b1110;
                    seg = 7'b0110001;
                end
            endcase
            if (!is_begin_manual_input && btnC_debouncer && !sorting) begin 
                is_begin_manual_input = 1;
            end else if (!sw[0] && !is_finished_manual_input) begin // Manual input mode 
                sorting <= 0;
                delay_counter <= 0;
                j <= 0;
                random_bars_generated <= 0; // Reset the flag
                sorted <= 0; // Reset the sorted flag
                if (!btnC && curr_index_manual < 5) begin 
                    curr_digit_manual = sw[9] ? 9 : sw[8] ? 8 : sw[7] ? 7 : sw[6] ? 6 : sw[5] ? 5 :
                                        sw[4] ? 4 : sw[3] ? 3 : sw[2] ? 2 : sw[1] ? 1 : 1;
                    bar_heights[curr_index_manual] <= curr_digit_manual * 7;
                    led[curr_index_manual] <= 1;
                end else if (btnC_debouncer) begin
                    led[curr_index_manual] <= 1;
                    curr_index_manual <= curr_index_manual + 1;
                    if (curr_index_manual == 5) 
                        is_finished_manual_input <= 1;
                end
            end else if (sw[0] && !btnL && !random_bars_generated) begin // Random input mode
                counter <= counter + 1; // Increment counter
                is_finished_manual_input = 0;
                for (i = 0; i < 5; i = i + 1) begin
                    bar_heights[i] <= (counter * 37 + i * 17) % 63 + 1; // Generate more random heights
                end
                sorting <= 0; // Ensure sorting is not started yet
                delay_counter <= 0;
                j <= 0;
                random_bars_generated <= 1; // Set the flag
                sorted <= 0; // Reset the sorted flag
            end else if (btnL && !sorting && !sorted && (is_finished_manual_input || random_bars_generated)) begin
                sorting <= 1; // Start sorting
                i <= 0; 
                j <= 0;
                dir <= 0;
            end else if (sorting) begin // Cocktail sort
                led[5:0] <= looping_leds; // Loading led
                if (looping_counter == 0) begin
                    looping_leds <= {looping_leds[3:0], looping_leds[4]};
                    looping_7_seg <= (looping_7_seg == 11) ? 0 : looping_7_seg + 1;
                end
                case (looping_7_seg) // Loading 7-seg
                    0: begin
                        an = 4'b0111;
                        seg = 7'b0111111;
                    end
                    1: begin
                        an = 4'b0111;
                        seg = 7'b1011111;
                    end
                    2: begin
                        an = 4'b0111;
                        seg = 7'b1101111;
                    end
                    3: begin
                        an = 4'b0111;
                        seg = 7'b1110111;
                    end
                    4: begin
                        an = 4'b1011;
                        seg = 7'b1110111;
                    end
                    5: begin
                        an = 4'b1101;
                        seg = 7'b1110111;
                    end
                    6: begin
                        an = 4'b1110;
                        seg = 7'b1110111;
                    end
                    7: begin
                        an = 4'b1110;
                        seg = 7'b1111011;
                    end
                    8: begin
                        an = 4'b1110;
                        seg = 7'b1111101;
                    end
                    9: begin
                        an = 4'b1110;
                        seg = 7'b0111111;
                    end
                    10: begin
                        an = 4'b1101;
                        seg = 7'b0111111;
                    end
                    11: begin
                        an = 4'b1011;
                        seg = 7'b0111111;
                    end
                endcase            
                if (delay_counter < SORT_DELAY) begin
                    delay_counter <= delay_counter + 1; // Increment delay counter
                end else begin
                    delay_counter <= 0; // Reset delay counter
                        if (dir == 0 && j < 4 - i) begin
                            if (bar_heights[j] > bar_heights[j + 1]) begin
                                // Swap adjacent bars if they are in the wrong order
                                {bar_heights[j], bar_heights[j + 1]} <= {bar_heights[j + 1], bar_heights[j]};
                                swap_from <= j;
                                swap_to <= j + 1; 
                                swap <= 1;
                            end else begin
                                swap_from <= 10;
                                swap_to <= 10; 
                                swap <= 0;                               
                            end
                            j <= j + 1; // Move to the next pair
                        end
                        else if (dir == 1 && j >= i - 1) begin 
                            if (bar_heights[j] > bar_heights[j + 1]) begin
                            // Swap adjacent bars if they are in the wrong order
                            {bar_heights[j], bar_heights[j + 1]} <= {bar_heights[j + 1], bar_heights[j]};
                            swap_from <= j;
                            swap_to <= j + 1; 
                            swap <= 1;
                        end else begin
                            swap_from <= 10;
                            swap_to <= 10; 
                            swap <= 0;                             
                        end
                        j <= j - 1; // Move to the next pair
                        end 
                    else begin
                        swap_from <= 10;
                        swap_to <= 10; 
                        swap <= 0;
                        if (i < 3) begin
                            //i <= i + 1; // Move to the next pass of the bubble sort
                            if (dir == 0) begin
                                j <= 3 - i; 
                                dir <= 1;
                                i <= i + 1;
                            end else begin
                                j <= 0;
                                dir <= 0;
                            end
                        end 
                        else begin
                            sorting <= 0; // Sorting is complete
                            sorted <= 1; // Set the sorted flag
                            is_finished_manual_input <= 0;
                            sorting_algorithm <= 4'b0011; // Display dOnE
                        end
                    end
                end
            end 
        end
        
        else if (sorting_algorithm == 4'b0011) begin // Done sorting
            case (anode_index)
                2'b00: begin
                    an = 4'b0111;
                    seg = 7'b0110000;
                end 
                2'b01: begin
                    an = 4'b1011;
                    seg = 7'b1101010;
                end
                2'b10: begin
                    an = 4'b1101;
                    seg = 7'b0000001;
                end 
                2'b11: begin
                    an = 4'b1110;
                    seg = 7'b1000010;
                end
            endcase
            led[5:0] <= 0;
        end 
        
        else if (sorting_algorithm == 4'b0000) begin // Start state
            case (anode_index) // Show Strt
                2'b00: begin
                    an = 4'b0111;
                    seg = 7'b1110000;
                end
                2'b01: begin
                    an = 4'b1011;
                    seg = 7'b1111010;
                end
                2'b10: begin
                    an = 4'b1101;
                    seg = 7'b1110000;
                end
                2'b11: begin
                    an = 4'b1110;
                    seg = 7'b0100100;
                end
            endcase
        end
    end
    
    //additional color definitions
    localparam YELLOW_COLOR = 16'hFFE0; // Yellow color
    localparam RED_COLOR = 16'hF800; // Red color
    localparam WHITE_COLOR = 16'hFFFF; // Red color
    integer bar_index;
    reg[6:0] vertical;
    reg [30:0] m_counter;
    reg [6:0] horizontal;
    integer TOTAL_MOVE;
    integer SPEED;
    
    //(m_counter == SORT_DELAY / (19 * (swap_to - swap_from)))
    always @(posedge clk) begin
    //params
    TOTAL_MOVE <= 19;
    SPEED <= 1_000_000;
    //
    if (sorting_algorithm == 4'b0010) begin
        TOTAL_MOVE <= 19 * (selection_sort_to - selection_sort_from);
    end
    if (delay_counter == 0) begin
        m_counter <= 0;
        movement <= 0;
    end
        if (swap == 1) begin
                m_counter <= m_counter + 1;
                if (m_counter == SPEED) begin
                    if (movement < TOTAL_MOVE) begin
                        movement <= movement + 1;
                    end

                    m_counter <= 0;
                end
            end
    end

    // Add more logic in the display block to change colors
    always @(*) begin
        horizontal = pixel_index % 96;
        vertical = pixel_index / 96;
        bar_index = ((pixel_index % 96) / (BAR_WIDTH + BAR_SPACING)) / 2;

        if (sorting_algorithm == 4'b0010) begin // selection sorting
            // First OLED
            if ((pixel_index % 96) < (BAR_WIDTH * 10 + BAR_SPACING * 9)) begin
                // Inside the bar area
                if (((pixel_index % 96) / (BAR_WIDTH + BAR_SPACING)) % 2 == 0) begin
                    if ((63 - (pixel_index / 96)) < bar_heights[((pixel_index % 96) / (BAR_WIDTH + BAR_SPACING)) / 2]) begin
                        if (sorting) begin
                            if ((((pixel_index % 96) / (BAR_WIDTH + BAR_SPACING)) / 2) == j - 1 && sorting) begin // If this is the selected bar, make it yellow
                                oled_data = YELLOW_COLOR;
                            end else if (((pixel_index % 96) / (BAR_WIDTH + BAR_SPACING)) / 2 < i) begin
                                oled_data = BAR_COLOR;
                            end else begin
                                oled_data = RED_COLOR;
                            end
                        end else begin
                            oled_data = BAR_COLOR;
                        end
                    end else begin
                        oled_data = BACKGROUND_COLOR;
                    end
                end else begin
                    oled_data = BACKGROUND_COLOR;
                end
            end else begin
                // Outside the bar area
                oled_data = BACKGROUND_COLOR;
            end    
        end
        else begin
            bar_index = ((pixel_index % 96) / (BAR_WIDTH + BAR_SPACING)) / 2; // Calculate the bar index
        
            // Default color is black(background)
            oled_data = BACKGROUND_COLOR;
            
            if ((pixel_index % 96) < (BAR_WIDTH * 10 + BAR_SPACING * 9)) begin // Inside the bar area
                if (((pixel_index % 96) / (BAR_WIDTH + BAR_SPACING)) % 2 == 0) begin // Inside a bar
                    if ((63 - (pixel_index / 96)) < bar_heights[bar_index]) begin
                        if (sorting_algorithm == 4'b0001) begin // bubble sorting
                            oled_data = BAR_COLOR;
                            // If sorting is in progress, color bars accordingly
                            if (sorting) begin
                                oled_data = RED_COLOR;
                                // If the bar is currently being compared, color it yellow
                                if (bar_index == j || bar_index == j + 1) begin
                                    oled_data = YELLOW_COLOR;
                                end
                                // If the bar is in the sorted position, color it red
                                if (bar_index >= 5 - i) begin
                                    oled_data = BAR_COLOR;
                                end
                            end
                        end
                        else if (sorting_algorithm == 4'b0100) begin //insertion sort
                            // Default bar color
                            oled_data = BAR_COLOR;
                            // If sorting is in progress, color bars accordingly
                            if (sorting) begin
                                oled_data = RED_COLOR; 
                                if (bar_index < i)
                                    oled_data = BAR_COLOR;   
                                if (bar_index == j || bar_index == j - 1)
                                    oled_data = YELLOW_COLOR;                             
                            end else if (sorted) begin
                                oled_data <= BAR_COLOR;
                            end
                            

                        end else if (sorting_algorithm == 4'b1000) begin //cocktail sort
                            oled_data = BAR_COLOR;
                            // If sorting is in progress, color bars accordingly
                            if (sorting) begin
                            //default sorting color = red
                                oled_data = RED_COLOR;
                                // If the bar is currently being compared, color it yellow
                                if (bar_index == j || bar_index == j + 1) begin
                                    oled_data = YELLOW_COLOR;
                                end
                
                                // If the bar is in the sorted position, color it red
                                if (bar_index >= 5 - i || bar_index < i && i==1 && dir == 0
                                || bar_index < i - 1 && i==2 && dir == 1
                                || bar_index < i && i==2 && dir == 0
                                || bar_index < i && i==3 && dir == 1
                                ) begin
                                    oled_data = BAR_COLOR;
                                end
                            end
                        end else if (sorting_algorithm == 4'b0011) begin //done sorting
                            if (sorted)
                                oled_data <= BAR_COLOR;
                        end
                    end
                end
            end
        end
        
    end
    
    
// 2nd OLED sorts, comment from here to debug so bitstream is faster
always @(*) begin
    if (sorting_algorithm == 0) begin
        // Your frame animation code goes here
            case (menuframe)
                0: begin
                    if (pixel_index2 == 97 || pixel_index2 == 99 || pixel_index2 == 101 || ((pixel_index2 >= 103) && (pixel_index2 <= 104)) || ((pixel_index2 >= 106) && (pixel_index2 <= 109)) || pixel_index2 == 111 || ((pixel_index2 >= 113) && (pixel_index2 <= 114)) || ((pixel_index2 >= 118) && (pixel_index2 <= 120)) || pixel_index2 == 195 || pixel_index2 == 197 || ((pixel_index2 >= 199) && (pixel_index2 <= 200)) || pixel_index2 == 202 || ((pixel_index2 >= 204) && (pixel_index2 <= 205)) || pixel_index2 == 207 || ((pixel_index2 >= 209) && (pixel_index2 <= 210)) || pixel_index2 == 213 || pixel_index2 == 289 || ((pixel_index2 >= 291) && (pixel_index2 <= 296)) || pixel_index2 == 298 || ((pixel_index2 >= 300) && (pixel_index2 <= 301)) || pixel_index2 == 303 || ((pixel_index2 >= 305) && (pixel_index2 <= 306)) || ((pixel_index2 >= 310) && (pixel_index2 <= 312)) || pixel_index2 == 385 || ((pixel_index2 >= 387) && (pixel_index2 <= 392)) || pixel_index2 == 394 || ((pixel_index2 >= 396) && (pixel_index2 <= 397)) || ((pixel_index2 >= 399) && (pixel_index2 <= 402)) || pixel_index2 == 408 || ((pixel_index2 >= 501) && (pixel_index2 <= 504)) || ((pixel_index2 >= 674) && (pixel_index2 <= 675)) || ((pixel_index2 >= 678) && (pixel_index2 <= 681)) || ((pixel_index2 >= 685) && (pixel_index2 <= 686)) || pixel_index2 == 688 || ((pixel_index2 >= 690) && (pixel_index2 <= 691)) || ((pixel_index2 >= 693) && (pixel_index2 <= 696)) || ((pixel_index2 >= 770) && (pixel_index2 <= 771)) || pixel_index2 == 774 || ((pixel_index2 >= 776) && (pixel_index2 <= 777)) || ((pixel_index2 >= 779) && (pixel_index2 <= 782)) || pixel_index2 == 784 || ((pixel_index2 >= 786) && (pixel_index2 <= 787)) || ((pixel_index2 >= 790) && (pixel_index2 <= 791)) || ((pixel_index2 >= 866) && (pixel_index2 <= 867)) || pixel_index2 == 870 || ((pixel_index2 >= 872) && (pixel_index2 <= 873)) || pixel_index2 == 875 || ((pixel_index2 >= 877) && (pixel_index2 <= 878)) || pixel_index2 == 880 || ((pixel_index2 >= 882) && (pixel_index2 <= 883)) || ((pixel_index2 >= 886) && (pixel_index2 <= 887)) || ((pixel_index2 >= 961) && (pixel_index2 <= 964)) || pixel_index2 == 966 || ((pixel_index2 >= 968) && (pixel_index2 <= 969)) || ((pixel_index2 >= 971) && (pixel_index2 <= 974)) || ((pixel_index2 >= 976) && (pixel_index2 <= 979)) || ((pixel_index2 >= 981) && (pixel_index2 <= 984)) || ((pixel_index2 >= 3938) && (pixel_index2 <= 3939)) || pixel_index2 == 3942 || pixel_index2 == 3945 || ((pixel_index2 >= 3947) && (pixel_index2 <= 3950)) || pixel_index2 == 3952 || ((pixel_index2 >= 3954) && (pixel_index2 <= 3955)) || ((pixel_index2 >= 3959) && (pixel_index2 <= 3962)) || ((pixel_index2 >= 3964) && (pixel_index2 <= 3967)) || ((pixel_index2 >= 3969) && (pixel_index2 <= 3972)) || ((pixel_index2 >= 3974) && (pixel_index2 <= 3977)) || pixel_index2 == 3979 || ((pixel_index2 >= 3981) && (pixel_index2 <= 3982)) || ((pixel_index2 >= 3984) && (pixel_index2 <= 3986)) || ((pixel_index2 >= 4034) && (pixel_index2 <= 4035)) || ((pixel_index2 >= 4039) && (pixel_index2 <= 4040)) || ((pixel_index2 >= 4045) && (pixel_index2 <= 4046)) || pixel_index2 == 4048 || ((pixel_index2 >= 4050) && (pixel_index2 <= 4051)) || ((pixel_index2 >= 4057) && (pixel_index2 <= 4058)) || ((pixel_index2 >= 4060) && (pixel_index2 <= 4061)) || pixel_index2 == 4065 || ((pixel_index2 >= 4067) && (pixel_index2 <= 4068)) || pixel_index2 == 4070 || ((pixel_index2 >= 4072) && (pixel_index2 <= 4073)) || ((pixel_index2 >= 4075) && (pixel_index2 <= 4078)) || ((pixel_index2 >= 4082) && (pixel_index2 <= 4083)) || ((pixel_index2 >= 4130) && (pixel_index2 <= 4131)) || ((pixel_index2 >= 4135) && (pixel_index2 <= 4136)) || ((pixel_index2 >= 4139) && (pixel_index2 <= 4140)) || pixel_index2 == 4142 || pixel_index2 == 4144 || ((pixel_index2 >= 4146) && (pixel_index2 <= 4147)) || ((pixel_index2 >= 4151) && (pixel_index2 <= 4152)) || pixel_index2 == 4154 || ((pixel_index2 >= 4157) && (pixel_index2 <= 4159)) || pixel_index2 == 4161 || ((pixel_index2 >= 4163) && (pixel_index2 <= 4164)) || pixel_index2 == 4166 || ((pixel_index2 >= 4168) && (pixel_index2 <= 4169)) || pixel_index2 == 4171 || ((pixel_index2 >= 4173) && (pixel_index2 <= 4174)) || ((pixel_index2 >= 4178) && (pixel_index2 <= 4179)) || ((pixel_index2 >= 4225) && (pixel_index2 <= 4228)) || pixel_index2 == 4230 || pixel_index2 == 4233 || ((pixel_index2 >= 4235) && (pixel_index2 <= 4238)) || ((pixel_index2 >= 4240) && (pixel_index2 <= 4243)) || ((pixel_index2 >= 4247) && (pixel_index2 <= 4250)) || ((pixel_index2 >= 4252) && (pixel_index2 <= 4254)) || ((pixel_index2 >= 4257) && (pixel_index2 <= 4260)) || ((pixel_index2 >= 4262) && (pixel_index2 <= 4265)) || pixel_index2 == 4267 || ((pixel_index2 >= 4269) && (pixel_index2 <= 4270)) || (pixel_index2 >= 4272) && (pixel_index2 <= 4274)) oled_data2 = 16'b1111001010010100;
                    else if (((pixel_index2 >= 124) && (pixel_index2 <= 190)) || ((pixel_index2 >= 220) && (pixel_index2 <= 221)) || pixel_index2 == 225 || pixel_index2 == 229 || pixel_index2 == 233 || pixel_index2 == 237 || pixel_index2 == 241 || pixel_index2 == 245 || pixel_index2 == 249 || pixel_index2 == 253 || pixel_index2 == 257 || pixel_index2 == 261 || pixel_index2 == 265 || pixel_index2 == 269 || pixel_index2 == 273 || pixel_index2 == 277 || pixel_index2 == 281 || ((pixel_index2 >= 285) && (pixel_index2 <= 286)) || ((pixel_index2 >= 316) && (pixel_index2 <= 317)) || pixel_index2 == 321 || pixel_index2 == 325 || pixel_index2 == 329 || pixel_index2 == 333 || pixel_index2 == 337 || pixel_index2 == 341 || pixel_index2 == 345 || pixel_index2 == 349 || pixel_index2 == 353 || pixel_index2 == 357 || pixel_index2 == 361 || pixel_index2 == 365 || pixel_index2 == 369 || pixel_index2 == 373 || pixel_index2 == 377 || ((pixel_index2 >= 381) && (pixel_index2 <= 382)) || ((pixel_index2 >= 412) && (pixel_index2 <= 413)) || pixel_index2 == 417 || pixel_index2 == 421 || pixel_index2 == 425 || pixel_index2 == 429 || pixel_index2 == 433 || pixel_index2 == 437 || pixel_index2 == 441 || pixel_index2 == 445 || pixel_index2 == 449 || pixel_index2 == 453 || pixel_index2 == 457 || pixel_index2 == 461 || pixel_index2 == 465 || pixel_index2 == 469 || pixel_index2 == 473 || ((pixel_index2 >= 477) && (pixel_index2 <= 478)) || ((pixel_index2 >= 508) && (pixel_index2 <= 509)) || pixel_index2 == 513 || pixel_index2 == 517 || pixel_index2 == 521 || pixel_index2 == 525 || pixel_index2 == 529 || pixel_index2 == 533 || pixel_index2 == 537 || pixel_index2 == 541 || pixel_index2 == 545 || pixel_index2 == 549 || pixel_index2 == 553 || pixel_index2 == 557 || pixel_index2 == 561 || pixel_index2 == 565 || pixel_index2 == 569 || ((pixel_index2 >= 573) && (pixel_index2 <= 574)) || ((pixel_index2 >= 604) && (pixel_index2 <= 605)) || pixel_index2 == 609 || pixel_index2 == 613 || pixel_index2 == 617 || pixel_index2 == 621 || pixel_index2 == 625 || pixel_index2 == 629 || pixel_index2 == 633 || pixel_index2 == 637 || pixel_index2 == 641 || pixel_index2 == 645 || pixel_index2 == 649 || pixel_index2 == 653 || pixel_index2 == 657 || pixel_index2 == 661 || pixel_index2 == 665 || ((pixel_index2 >= 669) && (pixel_index2 <= 670)) || ((pixel_index2 >= 700) && (pixel_index2 <= 701)) || pixel_index2 == 705 || pixel_index2 == 709 || pixel_index2 == 713 || pixel_index2 == 717 || pixel_index2 == 721 || pixel_index2 == 725 || pixel_index2 == 729 || pixel_index2 == 733 || pixel_index2 == 737 || pixel_index2 == 741 || pixel_index2 == 745 || pixel_index2 == 749 || pixel_index2 == 753 || pixel_index2 == 757 || pixel_index2 == 761 || ((pixel_index2 >= 765) && (pixel_index2 <= 766)) || ((pixel_index2 >= 796) && (pixel_index2 <= 862)) || ((pixel_index2 >= 892) && (pixel_index2 <= 894)) || ((pixel_index2 >= 897) && (pixel_index2 <= 898)) || ((pixel_index2 >= 901) && (pixel_index2 <= 902)) || ((pixel_index2 >= 905) && (pixel_index2 <= 906)) || ((pixel_index2 >= 909) && (pixel_index2 <= 910)) || ((pixel_index2 >= 913) && (pixel_index2 <= 914)) || ((pixel_index2 >= 917) && (pixel_index2 <= 918)) || ((pixel_index2 >= 921) && (pixel_index2 <= 922)) || ((pixel_index2 >= 925) && (pixel_index2 <= 926)) || ((pixel_index2 >= 929) && (pixel_index2 <= 930)) || ((pixel_index2 >= 933) && (pixel_index2 <= 934)) || ((pixel_index2 >= 937) && (pixel_index2 <= 938)) || ((pixel_index2 >= 941) && (pixel_index2 <= 942)) || ((pixel_index2 >= 945) && (pixel_index2 <= 946)) || ((pixel_index2 >= 949) && (pixel_index2 <= 950)) || ((pixel_index2 >= 953) && (pixel_index2 <= 954)) || ((pixel_index2 >= 957) && (pixel_index2 <= 958)) || ((pixel_index2 >= 988) && (pixel_index2 <= 1054)) || ((pixel_index2 >= 1084) && (pixel_index2 <= 1085)) || ((pixel_index2 >= 1087) && (pixel_index2 <= 1089)) || ((pixel_index2 >= 1091) && (pixel_index2 <= 1093)) || ((pixel_index2 >= 1095) && (pixel_index2 <= 1097)) || ((pixel_index2 >= 1099) && (pixel_index2 <= 1101)) || ((pixel_index2 >= 1103) && (pixel_index2 <= 1105)) || ((pixel_index2 >= 1107) && (pixel_index2 <= 1109)) || ((pixel_index2 >= 1111) && (pixel_index2 <= 1113)) || ((pixel_index2 >= 1115) && (pixel_index2 <= 1117)) || ((pixel_index2 >= 1119) && (pixel_index2 <= 1121)) || ((pixel_index2 >= 1123) && (pixel_index2 <= 1125)) || ((pixel_index2 >= 1127) && (pixel_index2 <= 1129)) || ((pixel_index2 >= 1131) && (pixel_index2 <= 1133)) || ((pixel_index2 >= 1135) && (pixel_index2 <= 1137)) || ((pixel_index2 >= 1139) && (pixel_index2 <= 1141)) || ((pixel_index2 >= 1143) && (pixel_index2 <= 1145)) || ((pixel_index2 >= 1147) && (pixel_index2 <= 1150)) || ((pixel_index2 >= 1182) && (pixel_index2 <= 1219)) || ((pixel_index2 >= 1240) && (pixel_index2 <= 1244)) || ((pixel_index2 >= 1278) && (pixel_index2 <= 1280)) || ((pixel_index2 >= 1283) && (pixel_index2 <= 1286)) || ((pixel_index2 >= 1290) && (pixel_index2 <= 1291)) || ((pixel_index2 >= 1293) && (pixel_index2 <= 1294)) || ((pixel_index2 >= 1314) && (pixel_index2 <= 1315)) || ((pixel_index2 >= 1336) && (pixel_index2 <= 1340)) || ((pixel_index2 >= 1374) && (pixel_index2 <= 1376)) || ((pixel_index2 >= 1378) && (pixel_index2 <= 1382)) || ((pixel_index2 >= 1386) && (pixel_index2 <= 1390)) || ((pixel_index2 >= 1410) && (pixel_index2 <= 1411)) || ((pixel_index2 >= 1432) && (pixel_index2 <= 1436)) || ((pixel_index2 >= 1470) && (pixel_index2 <= 1478)) || ((pixel_index2 >= 1482) && (pixel_index2 <= 1486)) || ((pixel_index2 >= 1506) && (pixel_index2 <= 1507)) || ((pixel_index2 >= 1528) && (pixel_index2 <= 1532)) || ((pixel_index2 >= 1566) && (pixel_index2 <= 1603)) || ((pixel_index2 >= 1624) && (pixel_index2 <= 1628)) || ((pixel_index2 >= 1662) && (pixel_index2 <= 1666)) || pixel_index2 == 1670 || pixel_index2 == 1674 || ((pixel_index2 >= 1678) && (pixel_index2 <= 1696)) || ((pixel_index2 >= 1698) && (pixel_index2 <= 1699)) || ((pixel_index2 >= 1720) && (pixel_index2 <= 1724)) || ((pixel_index2 >= 1758) && (pixel_index2 <= 1762)) || pixel_index2 == 1766 || pixel_index2 == 1770 || ((pixel_index2 >= 1774) && (pixel_index2 <= 1775)) || ((pixel_index2 >= 1777) && (pixel_index2 <= 1789)) || pixel_index2 == 1792 || ((pixel_index2 >= 1794) && (pixel_index2 <= 1795)) || pixel_index2 == 1816 || ((pixel_index2 >= 1818) && (pixel_index2 <= 1820)) || ((pixel_index2 >= 1854) && (pixel_index2 <= 1858)) || pixel_index2 == 1862 || pixel_index2 == 1866 || pixel_index2 == 1870 || ((pixel_index2 >= 1872) && (pixel_index2 <= 1878)) || ((pixel_index2 >= 1882) && (pixel_index2 <= 1888)) || ((pixel_index2 >= 1892) && (pixel_index2 <= 1913)) || ((pixel_index2 >= 1915) && (pixel_index2 <= 1916)) || ((pixel_index2 >= 1948) && (pixel_index2 <= 1973)) || pixel_index2 == 1988 || pixel_index2 == 1991 || ((pixel_index2 >= 1993) && (pixel_index2 <= 1994)) || pixel_index2 == 1996 || ((pixel_index2 >= 2000) && (pixel_index2 <= 2001)) || pixel_index2 == 2008 || ((pixel_index2 >= 2011) && (pixel_index2 <= 2014)) || ((pixel_index2 >= 2044) && (pixel_index2 <= 2046)) || ((pixel_index2 >= 2048) && (pixel_index2 <= 2054)) || ((pixel_index2 >= 2058) && (pixel_index2 <= 2069)) || ((pixel_index2 >= 2084) && (pixel_index2 <= 2085)) || pixel_index2 == 2089 || ((pixel_index2 >= 2091) && (pixel_index2 <= 2093)) || ((pixel_index2 >= 2095) && (pixel_index2 <= 2096)) || ((pixel_index2 >= 2104) && (pixel_index2 <= 2105)) || ((pixel_index2 >= 2107) && (pixel_index2 <= 2110)) || pixel_index2 == 2140 || pixel_index2 == 2142 || ((pixel_index2 >= 2144) && (pixel_index2 <= 2150)) || pixel_index2 == 2154 || ((pixel_index2 >= 2157) && (pixel_index2 <= 2168)) || pixel_index2 == 2178 || ((pixel_index2 >= 2180) && (pixel_index2 <= 2184)) || pixel_index2 == 2188 || ((pixel_index2 >= 2190) && (pixel_index2 <= 2192)) || ((pixel_index2 >= 2195) && (pixel_index2 <= 2197)) || ((pixel_index2 >= 2200) && (pixel_index2 <= 2206)) || ((pixel_index2 >= 2236) && (pixel_index2 <= 2238)) || ((pixel_index2 >= 2245) && (pixel_index2 <= 2246)) || pixel_index2 == 2250 || ((pixel_index2 >= 2252) && (pixel_index2 <= 2264)) || ((pixel_index2 >= 2274) && (pixel_index2 <= 2288)) || ((pixel_index2 >= 2291) && (pixel_index2 <= 2293)) || ((pixel_index2 >= 2296) && (pixel_index2 <= 2302)) || ((pixel_index2 >= 2332) && (pixel_index2 <= 2334)) || ((pixel_index2 >= 2341) && (pixel_index2 <= 2355)) || ((pixel_index2 >= 2374) && (pixel_index2 <= 2384)) || ((pixel_index2 >= 2392) && (pixel_index2 <= 2398)) || ((pixel_index2 >= 2428) && (pixel_index2 <= 2437)) || ((pixel_index2 >= 2443) && (pixel_index2 <= 2451)) || ((pixel_index2 >= 2470) && (pixel_index2 <= 2480)) || ((pixel_index2 >= 2487) && (pixel_index2 <= 2494)) || ((pixel_index2 >= 2526) && (pixel_index2 <= 2532)) || ((pixel_index2 >= 2540) && (pixel_index2 <= 2547)) || pixel_index2 == 2566 || ((pixel_index2 >= 2580) && (pixel_index2 <= 2588)) || ((pixel_index2 >= 2622) && (pixel_index2 <= 2626)) || pixel_index2 == 2636 || ((pixel_index2 >= 2639) && (pixel_index2 <= 2644)) || ((pixel_index2 >= 2647) && (pixel_index2 <= 2648)) || pixel_index2 == 2659 || ((pixel_index2 >= 2661) && (pixel_index2 <= 2662)) || ((pixel_index2 >= 2676) && (pixel_index2 <= 2684)) || ((pixel_index2 >= 2718) && (pixel_index2 <= 2721)) || pixel_index2 == 2732 || ((pixel_index2 >= 2735) && (pixel_index2 <= 2742)) || ((pixel_index2 >= 2756) && (pixel_index2 <= 2758)) || ((pixel_index2 >= 2772) && (pixel_index2 <= 2780)) || ((pixel_index2 >= 2814) && (pixel_index2 <= 2817)) || pixel_index2 == 2828 || ((pixel_index2 >= 2831) && (pixel_index2 <= 2838)) || ((pixel_index2 >= 2842) && (pixel_index2 <= 2848)) || ((pixel_index2 >= 2852) && (pixel_index2 <= 2859)) || ((pixel_index2 >= 2866) && (pixel_index2 <= 2876)) || ((pixel_index2 >= 2910) && (pixel_index2 <= 2913)) || pixel_index2 == 2924 || ((pixel_index2 >= 2927) && (pixel_index2 <= 2935)) || ((pixel_index2 >= 2938) && (pixel_index2 <= 2944)) || ((pixel_index2 >= 2947) && (pixel_index2 <= 2955)) || pixel_index2 == 2962 || ((pixel_index2 >= 2964) && (pixel_index2 <= 2972)) || ((pixel_index2 >= 3006) && (pixel_index2 <= 3013)) || ((pixel_index2 >= 3019) && (pixel_index2 <= 3021)) || ((pixel_index2 >= 3023) && (pixel_index2 <= 3032)) || ((pixel_index2 >= 3042) && (pixel_index2 <= 3051)) || ((pixel_index2 >= 3058) && (pixel_index2 <= 3060)) || pixel_index2 == 3063 || ((pixel_index2 >= 3065) && (pixel_index2 <= 3068)) || ((pixel_index2 >= 3102) && (pixel_index2 <= 3104)) || pixel_index2 == 3107 || ((pixel_index2 >= 3117) && (pixel_index2 <= 3123)) || ((pixel_index2 >= 3143) && (pixel_index2 <= 3147)) || ((pixel_index2 >= 3154) && (pixel_index2 <= 3155)) || pixel_index2 == 3159 || ((pixel_index2 >= 3161) && (pixel_index2 <= 3164)) || ((pixel_index2 >= 3198) && (pixel_index2 <= 3200)) || ((pixel_index2 >= 3202) && (pixel_index2 <= 3203)) || ((pixel_index2 >= 3213) && (pixel_index2 <= 3216)) || ((pixel_index2 >= 3218) && (pixel_index2 <= 3219)) || ((pixel_index2 >= 3239) && (pixel_index2 <= 3243)) || ((pixel_index2 >= 3250) && (pixel_index2 <= 3251)) || ((pixel_index2 >= 3255) && (pixel_index2 <= 3260)) || ((pixel_index2 >= 3292) && (pixel_index2 <= 3299)) || ((pixel_index2 >= 3309) && (pixel_index2 <= 3312)) || ((pixel_index2 >= 3314) && (pixel_index2 <= 3315)) || ((pixel_index2 >= 3335) && (pixel_index2 <= 3337)) || pixel_index2 == 3339 || ((pixel_index2 >= 3346) && (pixel_index2 <= 3347)) || ((pixel_index2 >= 3351) && (pixel_index2 <= 3352)) || ((pixel_index2 >= 3354) && (pixel_index2 <= 3358)) || ((pixel_index2 >= 3388) && (pixel_index2 <= 3393)) || pixel_index2 == 3395 || ((pixel_index2 >= 3405) && (pixel_index2 <= 3407)) || ((pixel_index2 >= 3409) && (pixel_index2 <= 3411)) || ((pixel_index2 >= 3431) && (pixel_index2 <= 3432)) || ((pixel_index2 >= 3434) && (pixel_index2 <= 3435)) || ((pixel_index2 >= 3438) && (pixel_index2 <= 3443)) || ((pixel_index2 >= 3447) && (pixel_index2 <= 3448)) || ((pixel_index2 >= 3450) && (pixel_index2 <= 3454)) || ((pixel_index2 >= 3484) && (pixel_index2 <= 3487)) || pixel_index2 == 3489 || pixel_index2 == 3491 || ((pixel_index2 >= 3501) && (pixel_index2 <= 3502)) || ((pixel_index2 >= 3505) && (pixel_index2 <= 3507)) || ((pixel_index2 >= 3527) && (pixel_index2 <= 3531)) || ((pixel_index2 >= 3538) && (pixel_index2 <= 3539)) || ((pixel_index2 >= 3543) && (pixel_index2 <= 3544)) || ((pixel_index2 >= 3546) && (pixel_index2 <= 3550)) || ((pixel_index2 >= 3580) && (pixel_index2 <= 3587)) || ((pixel_index2 >= 3597) && (pixel_index2 <= 3603)) || ((pixel_index2 >= 3623) && (pixel_index2 <= 3628)) || ((pixel_index2 >= 3633) && (pixel_index2 <= 3635)) || ((pixel_index2 >= 3639) && (pixel_index2 <= 3646)) || ((pixel_index2 >= 4620) && (pixel_index2 <= 4692)) || ((pixel_index2 >= 4707) && (pixel_index2 <= 4796)) || ((pixel_index2 >= 4803) && (pixel_index2 <= 4812)) || ((pixel_index2 >= 4814) && (pixel_index2 <= 4817)) || ((pixel_index2 >= 4819) && (pixel_index2 <= 4820)) || ((pixel_index2 >= 4827) && (pixel_index2 <= 4829)) || ((pixel_index2 >= 4834) && (pixel_index2 <= 4835)) || ((pixel_index2 >= 4838) && (pixel_index2 <= 4839)) || ((pixel_index2 >= 4841) && (pixel_index2 <= 4843)) || ((pixel_index2 >= 4845) && (pixel_index2 <= 4846)) || ((pixel_index2 >= 4851) && (pixel_index2 <= 4861)) || ((pixel_index2 >= 4863) && (pixel_index2 <= 4865)) || ((pixel_index2 >= 4868) && (pixel_index2 <= 4869)) || ((pixel_index2 >= 4871) && (pixel_index2 <= 4873)) || ((pixel_index2 >= 4880) && (pixel_index2 <= 4882)) || ((pixel_index2 >= 4887) && (pixel_index2 <= 4892)) || ((pixel_index2 >= 4899) && (pixel_index2 <= 4907)) || ((pixel_index2 >= 4910) && (pixel_index2 <= 4912)) || pixel_index2 == 4915 || pixel_index2 == 4924 || pixel_index2 == 4931 || pixel_index2 == 4935 || pixel_index2 == 4938 || pixel_index2 == 4941 || ((pixel_index2 >= 4948) && (pixel_index2 <= 4956)) || ((pixel_index2 >= 4959) && (pixel_index2 <= 4961)) || pixel_index2 == 4965 || pixel_index2 == 4968 || pixel_index2 == 4977 || ((pixel_index2 >= 4984) && (pixel_index2 <= 4988)) || ((pixel_index2 >= 4994) && (pixel_index2 <= 5003)) || ((pixel_index2 >= 5006) && (pixel_index2 <= 5008)) || pixel_index2 == 5011 || pixel_index2 == 5020 || pixel_index2 == 5027 || pixel_index2 == 5034 || pixel_index2 == 5037 || ((pixel_index2 >= 5044) && (pixel_index2 <= 5052)) || ((pixel_index2 >= 5055) && (pixel_index2 <= 5057)) || pixel_index2 == 5064 || pixel_index2 == 5073 || ((pixel_index2 >= 5080) && (pixel_index2 <= 5085)) || ((pixel_index2 >= 5090) && (pixel_index2 <= 5099)) || ((pixel_index2 >= 5102) && (pixel_index2 <= 5104)) || pixel_index2 == 5107 || ((pixel_index2 >= 5111) && (pixel_index2 <= 5112)) || ((pixel_index2 >= 5116) && (pixel_index2 <= 5119)) || ((pixel_index2 >= 5123) && (pixel_index2 <= 5124)) || pixel_index2 == 5130 || ((pixel_index2 >= 5133) && (pixel_index2 <= 5136)) || ((pixel_index2 >= 5140) && (pixel_index2 <= 5148)) || ((pixel_index2 >= 5151) && (pixel_index2 <= 5154)) || pixel_index2 == 5160 || ((pixel_index2 >= 5164) && (pixel_index2 <= 5165)) || pixel_index2 == 5169 || ((pixel_index2 >= 5173) && (pixel_index2 <= 5181)) || ((pixel_index2 >= 5186) && (pixel_index2 <= 5195)) || ((pixel_index2 >= 5198) && (pixel_index2 <= 5200)) || pixel_index2 == 5203 || ((pixel_index2 >= 5206) && (pixel_index2 <= 5209)) || ((pixel_index2 >= 5212) && (pixel_index2 <= 5216)) || ((pixel_index2 >= 5219) && (pixel_index2 <= 5220)) || pixel_index2 == 5226 || ((pixel_index2 >= 5229) && (pixel_index2 <= 5233)) || ((pixel_index2 >= 5236) && (pixel_index2 <= 5244)) || ((pixel_index2 >= 5247) && (pixel_index2 <= 5250)) || pixel_index2 == 5256 || ((pixel_index2 >= 5259) && (pixel_index2 <= 5262)) || pixel_index2 == 5265 || ((pixel_index2 >= 5271) && (pixel_index2 <= 5277)) || ((pixel_index2 >= 5282) && (pixel_index2 <= 5291)) || ((pixel_index2 >= 5294) && (pixel_index2 <= 5296)) || pixel_index2 == 5299 || ((pixel_index2 >= 5302) && (pixel_index2 <= 5305)) || ((pixel_index2 >= 5308) && (pixel_index2 <= 5312)) || pixel_index2 == 5315 || pixel_index2 == 5322 || ((pixel_index2 >= 5325) && (pixel_index2 <= 5329)) || ((pixel_index2 >= 5332) && (pixel_index2 <= 5340)) || ((pixel_index2 >= 5343) && (pixel_index2 <= 5345)) || pixel_index2 == 5352 || ((pixel_index2 >= 5355) && (pixel_index2 <= 5358)) || pixel_index2 == 5361 || ((pixel_index2 >= 5368) && (pixel_index2 <= 5373)) || ((pixel_index2 >= 5378) && (pixel_index2 <= 5387)) || ((pixel_index2 >= 5390) && (pixel_index2 <= 5392)) || pixel_index2 == 5395 || ((pixel_index2 >= 5398) && (pixel_index2 <= 5401)) || ((pixel_index2 >= 5404) && (pixel_index2 <= 5408)) || pixel_index2 == 5411 || pixel_index2 == 5415 || pixel_index2 == 5418 || ((pixel_index2 >= 5421) && (pixel_index2 <= 5425)) || ((pixel_index2 >= 5428) && (pixel_index2 <= 5436)) || ((pixel_index2 >= 5439) && (pixel_index2 <= 5441)) || pixel_index2 == 5445 || pixel_index2 == 5448 || ((pixel_index2 >= 5451) && (pixel_index2 <= 5454)) || ((pixel_index2 >= 5457) && (pixel_index2 <= 5458)) || ((pixel_index2 >= 5464) && (pixel_index2 <= 5469)) || ((pixel_index2 >= 5474) && (pixel_index2 <= 5483)) || ((pixel_index2 >= 5486) && (pixel_index2 <= 5488)) || pixel_index2 == 5491 || ((pixel_index2 >= 5494) && (pixel_index2 <= 5497)) || ((pixel_index2 >= 5500) && (pixel_index2 <= 5503)) || pixel_index2 == 5507 || ((pixel_index2 >= 5510) && (pixel_index2 <= 5511)) || pixel_index2 == 5514 || ((pixel_index2 >= 5517) && (pixel_index2 <= 5520)) || ((pixel_index2 >= 5524) && (pixel_index2 <= 5532)) || ((pixel_index2 >= 5535) && (pixel_index2 <= 5537)) || ((pixel_index2 >= 5540) && (pixel_index2 <= 5541)) || pixel_index2 == 5544 || ((pixel_index2 >= 5548) && (pixel_index2 <= 5549)) || ((pixel_index2 >= 5553) && (pixel_index2 <= 5556)) || ((pixel_index2 >= 5560) && (pixel_index2 <= 5565)) || ((pixel_index2 >= 5570) && (pixel_index2 <= 5575)) || pixel_index2 == 5584 || pixel_index2 == 5587 || ((pixel_index2 >= 5590) && (pixel_index2 <= 5593)) || pixel_index2 == 5596 || pixel_index2 == 5603 || pixel_index2 == 5610 || pixel_index2 == 5613 || ((pixel_index2 >= 5620) && (pixel_index2 <= 5624)) || pixel_index2 == 5633 || pixel_index2 == 5640 || pixel_index2 == 5649 || ((pixel_index2 >= 5656) && (pixel_index2 <= 5661)) || ((pixel_index2 >= 5667) && (pixel_index2 <= 5671)) || pixel_index2 == 5680 || pixel_index2 == 5683 || ((pixel_index2 >= 5686) && (pixel_index2 <= 5689)) || pixel_index2 == 5692 || pixel_index2 == 5699 || pixel_index2 == 5706 || pixel_index2 == 5709 || ((pixel_index2 >= 5716) && (pixel_index2 <= 5720)) || pixel_index2 == 5729 || pixel_index2 == 5736 || pixel_index2 == 5745 || ((pixel_index2 >= 5752) && (pixel_index2 <= 5756)) || ((pixel_index2 >= 5763) && (pixel_index2 <= 5768)) || ((pixel_index2 >= 5775) && (pixel_index2 <= 5776)) || ((pixel_index2 >= 5778) && (pixel_index2 <= 5780)) || ((pixel_index2 >= 5782) && (pixel_index2 <= 5785)) || ((pixel_index2 >= 5787) && (pixel_index2 <= 5789)) || ((pixel_index2 >= 5794) && (pixel_index2 <= 5796)) || ((pixel_index2 >= 5801) && (pixel_index2 <= 5802)) || ((pixel_index2 >= 5804) && (pixel_index2 <= 5806)) || ((pixel_index2 >= 5811) && (pixel_index2 <= 5817)) || ((pixel_index2 >= 5824) && (pixel_index2 <= 5826)) || ((pixel_index2 >= 5831) && (pixel_index2 <= 5833)) || ((pixel_index2 >= 5840) && (pixel_index2 <= 5842)) || ((pixel_index2 >= 5847) && (pixel_index2 <= 5852)) || (pixel_index2 >= 5868) && (pixel_index2 <= 5940)) oled_data2 = 16'b0000000000001010;
                    else if (pixel_index2 == 323 || pixel_index2 == 327 || pixel_index2 == 331 || pixel_index2 == 335 || pixel_index2 == 339 || pixel_index2 == 419 || pixel_index2 == 423 || pixel_index2 == 427 || pixel_index2 == 431 || pixel_index2 == 435 || pixel_index2 == 3253 || pixel_index2 == 3349) oled_data2 = 16'b0000010100000000;
                    else if (pixel_index2 == 511 || pixel_index2 == 535 || pixel_index2 == 539 || pixel_index2 == 543 || pixel_index2 == 547 || pixel_index2 == 551 || pixel_index2 == 555 || pixel_index2 == 559 || pixel_index2 == 563 || pixel_index2 == 567 || pixel_index2 == 571 || pixel_index2 == 607 || pixel_index2 == 631 || pixel_index2 == 635 || pixel_index2 == 639 || pixel_index2 == 643 || pixel_index2 == 647 || pixel_index2 == 651 || pixel_index2 == 655 || pixel_index2 == 659 || pixel_index2 == 663 || pixel_index2 == 667 || pixel_index2 == 3488) oled_data2 = 16'b1010000000000000;
                    else if (((pixel_index2 >= 895) && (pixel_index2 <= 896)) || ((pixel_index2 >= 899) && (pixel_index2 <= 900)) || ((pixel_index2 >= 903) && (pixel_index2 <= 904)) || ((pixel_index2 >= 907) && (pixel_index2 <= 908)) || ((pixel_index2 >= 911) && (pixel_index2 <= 912)) || ((pixel_index2 >= 915) && (pixel_index2 <= 916)) || ((pixel_index2 >= 919) && (pixel_index2 <= 920)) || ((pixel_index2 >= 923) && (pixel_index2 <= 924)) || ((pixel_index2 >= 927) && (pixel_index2 <= 928)) || ((pixel_index2 >= 931) && (pixel_index2 <= 932)) || ((pixel_index2 >= 935) && (pixel_index2 <= 936)) || ((pixel_index2 >= 939) && (pixel_index2 <= 940)) || ((pixel_index2 >= 943) && (pixel_index2 <= 944)) || ((pixel_index2 >= 947) && (pixel_index2 <= 948)) || ((pixel_index2 >= 951) && (pixel_index2 <= 952)) || ((pixel_index2 >= 955) && (pixel_index2 <= 956)) || ((pixel_index2 >= 3133) && (pixel_index2 <= 3134)) || pixel_index2 == 3228 || pixel_index2 == 3327 || ((pixel_index2 >= 3630) && (pixel_index2 <= 3631)) || pixel_index2 == 4802 || pixel_index2 == 4893 || pixel_index2 == 5762 || pixel_index2 == 5853) oled_data2 = 16'b1111011110011110;
                    else if (pixel_index2 == 1086 || pixel_index2 == 1287 || pixel_index2 == 1289 || pixel_index2 == 1479 || pixel_index2 == 1481 || pixel_index2 == 1667 || pixel_index2 == 1669 || pixel_index2 == 1671 || pixel_index2 == 1673 || pixel_index2 == 1675 || pixel_index2 == 1677 || pixel_index2 == 1859 || pixel_index2 == 1861 || pixel_index2 == 1863 || pixel_index2 == 1865 || pixel_index2 == 1867 || pixel_index2 == 1869 || ((pixel_index2 >= 1879) && (pixel_index2 <= 1881)) || ((pixel_index2 >= 1889) && (pixel_index2 <= 1891)) || ((pixel_index2 >= 1975) && (pixel_index2 <= 1987)) || ((pixel_index2 >= 2002) && (pixel_index2 <= 2007)) || pixel_index2 == 2055 || pixel_index2 == 2057 || ((pixel_index2 >= 2072) && (pixel_index2 <= 2073)) || ((pixel_index2 >= 2081) && (pixel_index2 <= 2082)) || ((pixel_index2 >= 2097) && (pixel_index2 <= 2103)) || pixel_index2 == 2169 || pixel_index2 == 2177 || ((pixel_index2 >= 2193) && (pixel_index2 <= 2194)) || ((pixel_index2 >= 2198) && (pixel_index2 <= 2199)) || pixel_index2 == 2239 || ((pixel_index2 >= 2241) && (pixel_index2 <= 2242)) || pixel_index2 == 2244 || pixel_index2 == 2247 || pixel_index2 == 2249 || pixel_index2 == 2265 || pixel_index2 == 2273 || ((pixel_index2 >= 2289) && (pixel_index2 <= 2290)) || ((pixel_index2 >= 2294) && (pixel_index2 <= 2295)) || pixel_index2 == 2335 || pixel_index2 == 2337 || pixel_index2 == 2339 || ((pixel_index2 >= 2356) && (pixel_index2 <= 2361)) || ((pixel_index2 >= 2369) && (pixel_index2 <= 2373)) || ((pixel_index2 >= 2385) && (pixel_index2 <= 2391)) || ((pixel_index2 >= 2438) && (pixel_index2 <= 2442)) || ((pixel_index2 >= 2452) && (pixel_index2 <= 2457)) || ((pixel_index2 >= 2465) && (pixel_index2 <= 2469)) || ((pixel_index2 >= 2481) && (pixel_index2 <= 2486)) || pixel_index2 == 2533 || pixel_index2 == 2539 || pixel_index2 == 2549 || ((pixel_index2 >= 2552) && (pixel_index2 <= 2553)) || pixel_index2 == 2561 || ((pixel_index2 >= 2564) && (pixel_index2 <= 2565)) || ((pixel_index2 >= 2627) && (pixel_index2 <= 2629)) || pixel_index2 == 2635 || ((pixel_index2 >= 2637) && (pixel_index2 <= 2638)) || pixel_index2 == 2649 || pixel_index2 == 2657 || ((pixel_index2 >= 2722) && (pixel_index2 <= 2725)) || pixel_index2 == 2731 || ((pixel_index2 >= 2733) && (pixel_index2 <= 2734)) || ((pixel_index2 >= 2743) && (pixel_index2 <= 2755)) || ((pixel_index2 >= 2818) && (pixel_index2 <= 2821)) || pixel_index2 == 2827 || ((pixel_index2 >= 2829) && (pixel_index2 <= 2830)) || ((pixel_index2 >= 2839) && (pixel_index2 <= 2841)) || ((pixel_index2 >= 2849) && (pixel_index2 <= 2851)) || ((pixel_index2 >= 2914) && (pixel_index2 <= 2917)) || pixel_index2 == 2923 || pixel_index2 == 2936 || pixel_index2 == 2945 || pixel_index2 == 2963 || ((pixel_index2 >= 3014) && (pixel_index2 <= 3018)) || ((pixel_index2 >= 3061) && (pixel_index2 <= 3062)) || pixel_index2 == 3064 || ((pixel_index2 >= 3108) && (pixel_index2 <= 3116)) || pixel_index2 == 3160 || ((pixel_index2 >= 3204) && (pixel_index2 <= 3212)) || ((pixel_index2 >= 3300) && (pixel_index2 <= 3308)) || pixel_index2 == 3317 || ((pixel_index2 >= 3319) && (pixel_index2 <= 3320)) || ((pixel_index2 >= 3330) && (pixel_index2 <= 3331)) || pixel_index2 == 3333 || pixel_index2 == 3338 || ((pixel_index2 >= 3396) && (pixel_index2 <= 3404)) || pixel_index2 == 3433 || ((pixel_index2 >= 3436) && (pixel_index2 <= 3437)) || ((pixel_index2 >= 3492) && (pixel_index2 <= 3500)) || ((pixel_index2 >= 3588) && (pixel_index2 <= 3596)) || ((pixel_index2 >= 3684) && (pixel_index2 <= 3692)) || ((pixel_index2 >= 3724) && (pixel_index2 <= 3729)) || ((pixel_index2 >= 3820) && (pixel_index2 <= 3825)) || ((pixel_index2 >= 3893) && (pixel_index2 <= 3894)) || ((pixel_index2 >= 3897) && (pixel_index2 <= 3905)) || ((pixel_index2 >= 3908) && (pixel_index2 <= 3909)) || ((pixel_index2 >= 3989) && (pixel_index2 <= 3990)) || ((pixel_index2 >= 3994) && (pixel_index2 <= 4000)) || ((pixel_index2 >= 4004) && (pixel_index2 <= 4005)) || ((pixel_index2 >= 4085) && (pixel_index2 <= 4086)) || ((pixel_index2 >= 4090) && (pixel_index2 <= 4096)) || ((pixel_index2 >= 4100) && (pixel_index2 <= 4101)) || pixel_index2 == 4706 || pixel_index2 == 4797 || pixel_index2 == 5666 || pixel_index2 == 5757) oled_data2 = 16'b0101001010001010;
                    else if (pixel_index2 == 1090 || pixel_index2 == 1094 || pixel_index2 == 1098 || pixel_index2 == 1102 || pixel_index2 == 1106) oled_data2 = 16'b1111011110001010;
                    else if (pixel_index2 == 1110 || pixel_index2 == 1114 || pixel_index2 == 1118 || pixel_index2 == 1122 || pixel_index2 == 1126 || pixel_index2 == 1130 || pixel_index2 == 1134 || pixel_index2 == 1138 || pixel_index2 == 1142 || pixel_index2 == 1146) oled_data2 = 16'b0000001010000000;
                    else if (pixel_index2 == 1155 || ((pixel_index2 >= 1159) && (pixel_index2 <= 1161)) || pixel_index2 == 1163 || ((pixel_index2 >= 1165) && (pixel_index2 <= 1166)) || pixel_index2 == 1168 || ((pixel_index2 >= 1170) && (pixel_index2 <= 1171)) || pixel_index2 == 1173 || ((pixel_index2 >= 1175) && (pixel_index2 <= 1176)) || pixel_index2 == 1254 || ((pixel_index2 >= 1256) && (pixel_index2 <= 1257)) || pixel_index2 == 1259 || ((pixel_index2 >= 1261) && (pixel_index2 <= 1262)) || ((pixel_index2 >= 1264) && (pixel_index2 <= 1267)) || ((pixel_index2 >= 1270) && (pixel_index2 <= 1272)) || pixel_index2 == 1350 || ((pixel_index2 >= 1352) && (pixel_index2 <= 1353)) || pixel_index2 == 1355 || ((pixel_index2 >= 1357) && (pixel_index2 <= 1358)) || pixel_index2 == 1360 || ((pixel_index2 >= 1362) && (pixel_index2 <= 1363)) || pixel_index2 == 1365 || ((pixel_index2 >= 1367) && (pixel_index2 <= 1368)) || ((pixel_index2 >= 1447) && (pixel_index2 <= 1449)) || ((pixel_index2 >= 1451) && (pixel_index2 <= 1454)) || ((pixel_index2 >= 1456) && (pixel_index2 <= 1459)) || (pixel_index2 >= 1461) && (pixel_index2 <= 1464)) oled_data2 = 16'b1010001010010100;
                    else if (((pixel_index2 >= 1281) && (pixel_index2 <= 1282)) || pixel_index2 == 1292 || pixel_index2 == 1295 || ((pixel_index2 >= 1297) && (pixel_index2 <= 1299)) || pixel_index2 == 1302 || ((pixel_index2 >= 1304) && (pixel_index2 <= 1305)) || pixel_index2 == 1307 || pixel_index2 == 1309 || pixel_index2 == 1311 || pixel_index2 == 1313 || pixel_index2 == 1377 || ((pixel_index2 >= 1392) && (pixel_index2 <= 1395)) || ((pixel_index2 >= 1397) && (pixel_index2 <= 1399)) || pixel_index2 == 1401 || ((pixel_index2 >= 1403) && (pixel_index2 <= 1404)) || pixel_index2 == 1406 || pixel_index2 == 1409 || ((pixel_index2 >= 1487) && (pixel_index2 <= 1488)) || pixel_index2 == 1490 || pixel_index2 == 1493 || pixel_index2 == 1495 || pixel_index2 == 1497 || ((pixel_index2 >= 1499) && (pixel_index2 <= 1500)) || ((pixel_index2 >= 1502) && (pixel_index2 <= 1503)) || pixel_index2 == 1505 || pixel_index2 == 1697 || pixel_index2 == 1776 || ((pixel_index2 >= 1790) && (pixel_index2 <= 1791)) || pixel_index2 == 1793 || pixel_index2 == 1817 || pixel_index2 == 1871 || pixel_index2 == 1914 || pixel_index2 == 1974 || ((pixel_index2 >= 1989) && (pixel_index2 <= 1990)) || pixel_index2 == 1992 || pixel_index2 == 1995 || ((pixel_index2 >= 1997) && (pixel_index2 <= 1999)) || ((pixel_index2 >= 2009) && (pixel_index2 <= 2010)) || pixel_index2 == 2047 || ((pixel_index2 >= 2070) && (pixel_index2 <= 2071)) || pixel_index2 == 2083 || ((pixel_index2 >= 2086) && (pixel_index2 <= 2088)) || pixel_index2 == 2090 || pixel_index2 == 2094 || pixel_index2 == 2106 || pixel_index2 == 2141 || pixel_index2 == 2143 || ((pixel_index2 >= 2155) && (pixel_index2 <= 2156)) || pixel_index2 == 2179 || ((pixel_index2 >= 2185) && (pixel_index2 <= 2187)) || pixel_index2 == 2189 || pixel_index2 == 2240 || pixel_index2 == 2243 || pixel_index2 == 2251 || pixel_index2 == 2336 || pixel_index2 == 2338 || pixel_index2 == 2340 || pixel_index2 == 2548 || ((pixel_index2 >= 2550) && (pixel_index2 <= 2551)) || ((pixel_index2 >= 2562) && (pixel_index2 <= 2563)) || ((pixel_index2 >= 2567) && (pixel_index2 <= 2579)) || ((pixel_index2 >= 2645) && (pixel_index2 <= 2646)) || pixel_index2 == 2658 || pixel_index2 == 2660 || ((pixel_index2 >= 2663) && (pixel_index2 <= 2675)) || ((pixel_index2 >= 2759) && (pixel_index2 <= 2771)) || ((pixel_index2 >= 2925) && (pixel_index2 <= 2926)) || pixel_index2 == 2937 || pixel_index2 == 2946 || pixel_index2 == 3022 || ((pixel_index2 >= 3105) && (pixel_index2 <= 3106)) || pixel_index2 == 3201 || pixel_index2 == 3217 || ((pixel_index2 >= 3230) && (pixel_index2 <= 3231)) || pixel_index2 == 3313 || pixel_index2 == 3324 || pixel_index2 == 3408 || ((pixel_index2 >= 3421) && (pixel_index2 <= 3422)) || ((pixel_index2 >= 3503) && (pixel_index2 <= 3504)) || ((pixel_index2 >= 3533) && (pixel_index2 <= 3536)) || pixel_index2 == 3629 || pixel_index2 == 3632) oled_data2 = 16'b1010010100010100;
                    else if (pixel_index2 == 1296 || ((pixel_index2 >= 1300) && (pixel_index2 <= 1301)) || pixel_index2 == 1303 || pixel_index2 == 1306 || pixel_index2 == 1308 || pixel_index2 == 1310 || pixel_index2 == 1312 || pixel_index2 == 1391 || pixel_index2 == 1396 || pixel_index2 == 1400 || pixel_index2 == 1402 || pixel_index2 == 1405 || ((pixel_index2 >= 1407) && (pixel_index2 <= 1408)) || pixel_index2 == 1489 || ((pixel_index2 >= 1491) && (pixel_index2 <= 1492)) || pixel_index2 == 1494 || pixel_index2 == 1496 || pixel_index2 == 1498 || pixel_index2 == 1501 || pixel_index2 == 1504 || pixel_index2 == 3353 || pixel_index2 == 3449 || pixel_index2 == 3545) oled_data2 = 16'b0101001010010100;
                    else if (((pixel_index2 >= 1317) && (pixel_index2 <= 1319)) || pixel_index2 == 1324 || ((pixel_index2 >= 1327) && (pixel_index2 <= 1329)) || ((pixel_index2 >= 1332) && (pixel_index2 <= 1334)) || pixel_index2 == 1415 || pixel_index2 == 1420 || pixel_index2 == 1425 || pixel_index2 == 1428 || ((pixel_index2 >= 1509) && (pixel_index2 <= 1511)) || ((pixel_index2 >= 1514) && (pixel_index2 <= 1516)) || ((pixel_index2 >= 1519) && (pixel_index2 <= 1521)) || ((pixel_index2 >= 1524) && (pixel_index2 <= 1526)) || pixel_index2 == 1607 || pixel_index2 == 1617 || pixel_index2 == 1622 || pixel_index2 == 1703 || pixel_index2 == 1713 || (pixel_index2 >= 1716) && (pixel_index2 <= 1718)) oled_data2 = 16'b1010000000001010;
                    else if (((pixel_index2 >= 1637) && (pixel_index2 <= 1638)) || ((pixel_index2 >= 1641) && (pixel_index2 <= 1644)) || ((pixel_index2 >= 1646) && (pixel_index2 <= 1649)) || ((pixel_index2 >= 1652) && (pixel_index2 <= 1654)) || pixel_index2 == 1732 || pixel_index2 == 1735 || pixel_index2 == 1740 || pixel_index2 == 1745 || pixel_index2 == 1747 || pixel_index2 == 1831 || pixel_index2 == 1836 || ((pixel_index2 >= 1839) && (pixel_index2 <= 1841)) || ((pixel_index2 >= 1844) && (pixel_index2 <= 1845)) || pixel_index2 == 1924 || pixel_index2 == 1927 || pixel_index2 == 1932 || pixel_index2 == 1937 || pixel_index2 == 1942 || ((pixel_index2 >= 2021) && (pixel_index2 <= 2022)) || pixel_index2 == 2028 || ((pixel_index2 >= 2030) && (pixel_index2 <= 2033)) || (pixel_index2 >= 2035) && (pixel_index2 <= 2037)) oled_data2 = 16'b0101010100011110;
                    else if (pixel_index2 == 2213 || pixel_index2 == 2216 || ((pixel_index2 >= 2219) && (pixel_index2 <= 2221)) || pixel_index2 == 2223 || pixel_index2 == 2226 || ((pixel_index2 >= 2228) && (pixel_index2 <= 2230)) || pixel_index2 == 2310 || pixel_index2 == 2312 || pixel_index2 == 2314 || pixel_index2 == 2319 || pixel_index2 == 2322 || pixel_index2 == 2325 || ((pixel_index2 >= 2406) && (pixel_index2 <= 2408)) || ((pixel_index2 >= 2411) && (pixel_index2 <= 2412)) || ((pixel_index2 >= 2415) && (pixel_index2 <= 2416)) || pixel_index2 == 2418 || pixel_index2 == 2421 || pixel_index2 == 2501 || pixel_index2 == 2504 || pixel_index2 == 2509 || pixel_index2 == 2511 || ((pixel_index2 >= 2513) && (pixel_index2 <= 2514)) || pixel_index2 == 2517 || ((pixel_index2 >= 2598) && (pixel_index2 <= 2600)) || ((pixel_index2 >= 2602) && (pixel_index2 <= 2604)) || pixel_index2 == 2607 || pixel_index2 == 2610 || (pixel_index2 >= 2612) && (pixel_index2 <= 2614)) oled_data2 = 16'b1010011110001010;
                    else if (pixel_index2 == 2788 || pixel_index2 == 2791 || ((pixel_index2 >= 2794) && (pixel_index2 <= 2795)) || ((pixel_index2 >= 2799) && (pixel_index2 <= 2800)) || ((pixel_index2 >= 2804) && (pixel_index2 <= 2805)) || pixel_index2 == 2885 || pixel_index2 == 2887 || pixel_index2 == 2889 || pixel_index2 == 2892 || pixel_index2 == 2894 || pixel_index2 == 2897 || pixel_index2 == 2899 || pixel_index2 == 2902 || ((pixel_index2 >= 2982) && (pixel_index2 <= 2983)) || pixel_index2 == 2988 || pixel_index2 == 2990 || pixel_index2 == 2993 || pixel_index2 == 2998 || pixel_index2 == 3077 || pixel_index2 == 3079 || pixel_index2 == 3081 || pixel_index2 == 3084 || pixel_index2 == 3086 || pixel_index2 == 3089 || pixel_index2 == 3091 || pixel_index2 == 3094 || pixel_index2 == 3172 || pixel_index2 == 3175 || ((pixel_index2 >= 3178) && (pixel_index2 <= 3179)) || ((pixel_index2 >= 3183) && (pixel_index2 <= 3184)) || (pixel_index2 >= 3188) && (pixel_index2 <= 3189)) oled_data2 = 16'b1111010100001010;
                    else if (pixel_index2 == 3229 || (pixel_index2 >= 3325) && (pixel_index2 <= 3326)) oled_data2 = 16'b0101010100001010;
                    else if (((pixel_index2 >= 3364) && (pixel_index2 <= 3367)) || ((pixel_index2 >= 3370) && (pixel_index2 <= 3372)) || ((pixel_index2 >= 3375) && (pixel_index2 <= 3376)) || ((pixel_index2 >= 3380) && (pixel_index2 <= 3382)) || pixel_index2 == 3463 || pixel_index2 == 3465 || pixel_index2 == 3468 || pixel_index2 == 3470 || pixel_index2 == 3473 || pixel_index2 == 3475 || pixel_index2 == 3478 || pixel_index2 == 3559 || ((pixel_index2 >= 3562) && (pixel_index2 <= 3564)) || pixel_index2 == 3566 || pixel_index2 == 3569 || ((pixel_index2 >= 3572) && (pixel_index2 <= 3574)) || pixel_index2 == 3655 || pixel_index2 == 3657 || pixel_index2 == 3660 || pixel_index2 == 3662 || pixel_index2 == 3665 || pixel_index2 == 3667 || pixel_index2 == 3670 || pixel_index2 == 3751 || ((pixel_index2 >= 3754) && (pixel_index2 <= 3756)) || pixel_index2 == 3758 || pixel_index2 == 3761 || (pixel_index2 >= 3764) && (pixel_index2 <= 3766)) oled_data2 = 16'b1010001010001010;
                    else if (pixel_index2 == 3394 || pixel_index2 == 3490) oled_data2 = 16'b0000000000010100;
                    else if (pixel_index2 == 3532 || pixel_index2 == 3537) oled_data2 = 16'b0101000000000000;
                    else if (((pixel_index2 >= 4008) && (pixel_index2 <= 4009)) || ((pixel_index2 >= 4012) && (pixel_index2 <= 4015)) || ((pixel_index2 >= 4017) && (pixel_index2 <= 4020)) || ((pixel_index2 >= 4022) && (pixel_index2 <= 4025)) || pixel_index2 == 4027 || ((pixel_index2 >= 4029) && (pixel_index2 <= 4030)) || ((pixel_index2 >= 4104) && (pixel_index2 <= 4105)) || ((pixel_index2 >= 4110) && (pixel_index2 <= 4111)) || ((pixel_index2 >= 4113) && (pixel_index2 <= 4114)) || ((pixel_index2 >= 4120) && (pixel_index2 <= 4121)) || ((pixel_index2 >= 4124) && (pixel_index2 <= 4126)) || ((pixel_index2 >= 4200) && (pixel_index2 <= 4201)) || ((pixel_index2 >= 4204) && (pixel_index2 <= 4205)) || pixel_index2 == 4207 || ((pixel_index2 >= 4210) && (pixel_index2 <= 4212)) || ((pixel_index2 >= 4214) && (pixel_index2 <= 4215)) || pixel_index2 == 4217 || pixel_index2 == 4219 || ((pixel_index2 >= 4221) && (pixel_index2 <= 4222)) || ((pixel_index2 >= 4295) && (pixel_index2 <= 4298)) || ((pixel_index2 >= 4300) && (pixel_index2 <= 4303)) || ((pixel_index2 >= 4305) && (pixel_index2 <= 4307)) || ((pixel_index2 >= 4310) && (pixel_index2 <= 4313)) || (pixel_index2 >= 4315) && (pixel_index2 <= 4318)) oled_data2 = 16'b0101011110010100;
                    else if (((pixel_index2 >= 4423) && (pixel_index2 <= 4505)) || ((pixel_index2 >= 4513) && (pixel_index2 <= 4518)) || (pixel_index2 >= 4602) && (pixel_index2 <= 4606)) oled_data2 = 16'b0000001010011110;
                    else if (((pixel_index2 >= 4519) && (pixel_index2 <= 4601)) || ((pixel_index2 >= 4609) && (pixel_index2 <= 4619)) || ((pixel_index2 >= 4693) && (pixel_index2 <= 4702)) || pixel_index2 == 4705 || pixel_index2 == 4798 || pixel_index2 == 4801 || pixel_index2 == 4894 || ((pixel_index2 >= 4897) && (pixel_index2 <= 4898)) || ((pixel_index2 >= 4989) && (pixel_index2 <= 4990)) || pixel_index2 == 4993 || pixel_index2 == 5086 || pixel_index2 == 5089 || pixel_index2 == 5182 || pixel_index2 == 5185 || pixel_index2 == 5278 || pixel_index2 == 5281 || pixel_index2 == 5374 || pixel_index2 == 5377 || pixel_index2 == 5470 || pixel_index2 == 5473 || pixel_index2 == 5566 || pixel_index2 == 5569 || pixel_index2 == 5662 || pixel_index2 == 5665 || pixel_index2 == 5758 || pixel_index2 == 5761 || pixel_index2 == 5854 || ((pixel_index2 >= 5857) && (pixel_index2 <= 5867)) || ((pixel_index2 >= 5941) && (pixel_index2 <= 5950)) || (pixel_index2 >= 5959) && (pixel_index2 <= 6041)) oled_data2 = 16'b0000001010010100;
                    else if (pixel_index2 == 4813 || pixel_index2 == 4818 || ((pixel_index2 >= 4821) && (pixel_index2 <= 4826)) || ((pixel_index2 >= 4830) && (pixel_index2 <= 4833)) || ((pixel_index2 >= 4836) && (pixel_index2 <= 4837)) || pixel_index2 == 4840 || pixel_index2 == 4844 || ((pixel_index2 >= 4847) && (pixel_index2 <= 4850)) || pixel_index2 == 4862 || ((pixel_index2 >= 4866) && (pixel_index2 <= 4867)) || pixel_index2 == 4870 || ((pixel_index2 >= 4874) && (pixel_index2 <= 4879)) || ((pixel_index2 >= 4883) && (pixel_index2 <= 4886)) || pixel_index2 == 4908 || pixel_index2 == 4913 || pixel_index2 == 4916 || pixel_index2 == 4923 || pixel_index2 == 4925 || pixel_index2 == 4930 || pixel_index2 == 4934 || pixel_index2 == 4937 || pixel_index2 == 4939 || pixel_index2 == 4942 || pixel_index2 == 4947 || pixel_index2 == 4957 || pixel_index2 == 4964 || pixel_index2 == 4967 || pixel_index2 == 4969 || pixel_index2 == 4976 || pixel_index2 == 4978 || pixel_index2 == 4983 || pixel_index2 == 5031 || pixel_index2 == 5061 || pixel_index2 == 5221 || pixel_index2 == 5251 || ((pixel_index2 >= 5268) && (pixel_index2 <= 5270)) || pixel_index2 == 5316 || pixel_index2 == 5346 || pixel_index2 == 5367 || pixel_index2 == 5504 || pixel_index2 == 5521 || pixel_index2 == 5547 || pixel_index2 == 5550 || pixel_index2 == 5557 || ((pixel_index2 >= 5576) && (pixel_index2 <= 5579)) || ((pixel_index2 >= 5582) && (pixel_index2 <= 5583)) || ((pixel_index2 >= 5597) && (pixel_index2 <= 5599)) || ((pixel_index2 >= 5606) && (pixel_index2 <= 5607)) || ((pixel_index2 >= 5614) && (pixel_index2 <= 5616)) || ((pixel_index2 >= 5625) && (pixel_index2 <= 5628)) || ((pixel_index2 >= 5631) && (pixel_index2 <= 5632)) || ((pixel_index2 >= 5636) && (pixel_index2 <= 5637)) || ((pixel_index2 >= 5644) && (pixel_index2 <= 5645)) || (pixel_index2 >= 5650) && (pixel_index2 <= 5652)) oled_data2 = 16'b0101001010000000;
                    else if (pixel_index2 == 4909 || pixel_index2 == 4914 || ((pixel_index2 >= 4917) && (pixel_index2 <= 4922)) || ((pixel_index2 >= 4926) && (pixel_index2 <= 4929)) || ((pixel_index2 >= 4932) && (pixel_index2 <= 4933)) || pixel_index2 == 4936 || pixel_index2 == 4940 || ((pixel_index2 >= 4943) && (pixel_index2 <= 4946)) || pixel_index2 == 4958 || ((pixel_index2 >= 4962) && (pixel_index2 <= 4963)) || pixel_index2 == 4966 || ((pixel_index2 >= 4970) && (pixel_index2 <= 4975)) || ((pixel_index2 >= 4979) && (pixel_index2 <= 4982)) || ((pixel_index2 >= 5004) && (pixel_index2 <= 5005)) || ((pixel_index2 >= 5009) && (pixel_index2 <= 5010)) || ((pixel_index2 >= 5012) && (pixel_index2 <= 5019)) || ((pixel_index2 >= 5021) && (pixel_index2 <= 5026)) || ((pixel_index2 >= 5028) && (pixel_index2 <= 5030)) || ((pixel_index2 >= 5032) && (pixel_index2 <= 5033)) || ((pixel_index2 >= 5035) && (pixel_index2 <= 5036)) || ((pixel_index2 >= 5038) && (pixel_index2 <= 5043)) || ((pixel_index2 >= 5053) && (pixel_index2 <= 5054)) || ((pixel_index2 >= 5058) && (pixel_index2 <= 5060)) || ((pixel_index2 >= 5062) && (pixel_index2 <= 5063)) || ((pixel_index2 >= 5065) && (pixel_index2 <= 5072)) || ((pixel_index2 >= 5074) && (pixel_index2 <= 5079)) || ((pixel_index2 >= 5100) && (pixel_index2 <= 5101)) || ((pixel_index2 >= 5105) && (pixel_index2 <= 5106)) || ((pixel_index2 >= 5108) && (pixel_index2 <= 5110)) || ((pixel_index2 >= 5113) && (pixel_index2 <= 5115)) || ((pixel_index2 >= 5120) && (pixel_index2 <= 5122)) || ((pixel_index2 >= 5125) && (pixel_index2 <= 5129)) || ((pixel_index2 >= 5131) && (pixel_index2 <= 5132)) || ((pixel_index2 >= 5137) && (pixel_index2 <= 5139)) || ((pixel_index2 >= 5149) && (pixel_index2 <= 5150)) || ((pixel_index2 >= 5155) && (pixel_index2 <= 5159)) || ((pixel_index2 >= 5161) && (pixel_index2 <= 5163)) || ((pixel_index2 >= 5166) && (pixel_index2 <= 5168)) || ((pixel_index2 >= 5170) && (pixel_index2 <= 5172)) || ((pixel_index2 >= 5196) && (pixel_index2 <= 5197)) || ((pixel_index2 >= 5201) && (pixel_index2 <= 5202)) || ((pixel_index2 >= 5204) && (pixel_index2 <= 5205)) || ((pixel_index2 >= 5210) && (pixel_index2 <= 5211)) || ((pixel_index2 >= 5217) && (pixel_index2 <= 5218)) || ((pixel_index2 >= 5222) && (pixel_index2 <= 5225)) || ((pixel_index2 >= 5227) && (pixel_index2 <= 5228)) || ((pixel_index2 >= 5234) && (pixel_index2 <= 5235)) || ((pixel_index2 >= 5245) && (pixel_index2 <= 5246)) || ((pixel_index2 >= 5252) && (pixel_index2 <= 5255)) || ((pixel_index2 >= 5257) && (pixel_index2 <= 5258)) || ((pixel_index2 >= 5263) && (pixel_index2 <= 5264)) || ((pixel_index2 >= 5266) && (pixel_index2 <= 5267)) || ((pixel_index2 >= 5292) && (pixel_index2 <= 5293)) || ((pixel_index2 >= 5297) && (pixel_index2 <= 5298)) || ((pixel_index2 >= 5300) && (pixel_index2 <= 5301)) || ((pixel_index2 >= 5306) && (pixel_index2 <= 5307)) || ((pixel_index2 >= 5313) && (pixel_index2 <= 5314)) || ((pixel_index2 >= 5317) && (pixel_index2 <= 5321)) || ((pixel_index2 >= 5323) && (pixel_index2 <= 5324)) || ((pixel_index2 >= 5330) && (pixel_index2 <= 5331)) || ((pixel_index2 >= 5341) && (pixel_index2 <= 5342)) || ((pixel_index2 >= 5347) && (pixel_index2 <= 5351)) || ((pixel_index2 >= 5353) && (pixel_index2 <= 5354)) || ((pixel_index2 >= 5359) && (pixel_index2 <= 5360)) || ((pixel_index2 >= 5362) && (pixel_index2 <= 5366)) || ((pixel_index2 >= 5388) && (pixel_index2 <= 5389)) || ((pixel_index2 >= 5393) && (pixel_index2 <= 5394)) || ((pixel_index2 >= 5396) && (pixel_index2 <= 5397)) || ((pixel_index2 >= 5402) && (pixel_index2 <= 5403)) || ((pixel_index2 >= 5409) && (pixel_index2 <= 5410)) || ((pixel_index2 >= 5412) && (pixel_index2 <= 5414)) || ((pixel_index2 >= 5416) && (pixel_index2 <= 5417)) || ((pixel_index2 >= 5419) && (pixel_index2 <= 5420)) || ((pixel_index2 >= 5426) && (pixel_index2 <= 5427)) || ((pixel_index2 >= 5437) && (pixel_index2 <= 5438)) || ((pixel_index2 >= 5442) && (pixel_index2 <= 5444)) || ((pixel_index2 >= 5446) && (pixel_index2 <= 5447)) || ((pixel_index2 >= 5449) && (pixel_index2 <= 5450)) || ((pixel_index2 >= 5455) && (pixel_index2 <= 5456)) || ((pixel_index2 >= 5459) && (pixel_index2 <= 5463)) || ((pixel_index2 >= 5484) && (pixel_index2 <= 5485)) || ((pixel_index2 >= 5489) && (pixel_index2 <= 5490)) || ((pixel_index2 >= 5492) && (pixel_index2 <= 5493)) || ((pixel_index2 >= 5498) && (pixel_index2 <= 5499)) || ((pixel_index2 >= 5505) && (pixel_index2 <= 5506)) || ((pixel_index2 >= 5508) && (pixel_index2 <= 5509)) || ((pixel_index2 >= 5512) && (pixel_index2 <= 5513)) || ((pixel_index2 >= 5515) && (pixel_index2 <= 5516)) || ((pixel_index2 >= 5522) && (pixel_index2 <= 5523)) || ((pixel_index2 >= 5533) && (pixel_index2 <= 5534)) || ((pixel_index2 >= 5538) && (pixel_index2 <= 5539)) || ((pixel_index2 >= 5542) && (pixel_index2 <= 5543)) || ((pixel_index2 >= 5545) && (pixel_index2 <= 5546)) || ((pixel_index2 >= 5551) && (pixel_index2 <= 5552)) || ((pixel_index2 >= 5558) && (pixel_index2 <= 5559)) || ((pixel_index2 >= 5580) && (pixel_index2 <= 5581)) || ((pixel_index2 >= 5585) && (pixel_index2 <= 5586)) || ((pixel_index2 >= 5588) && (pixel_index2 <= 5589)) || ((pixel_index2 >= 5594) && (pixel_index2 <= 5595)) || ((pixel_index2 >= 5600) && (pixel_index2 <= 5602)) || ((pixel_index2 >= 5604) && (pixel_index2 <= 5605)) || ((pixel_index2 >= 5608) && (pixel_index2 <= 5609)) || ((pixel_index2 >= 5611) && (pixel_index2 <= 5612)) || ((pixel_index2 >= 5617) && (pixel_index2 <= 5619)) || ((pixel_index2 >= 5629) && (pixel_index2 <= 5630)) || ((pixel_index2 >= 5634) && (pixel_index2 <= 5635)) || ((pixel_index2 >= 5638) && (pixel_index2 <= 5639)) || ((pixel_index2 >= 5641) && (pixel_index2 <= 5643)) || ((pixel_index2 >= 5646) && (pixel_index2 <= 5648)) || ((pixel_index2 >= 5653) && (pixel_index2 <= 5655)) || ((pixel_index2 >= 5672) && (pixel_index2 <= 5679)) || ((pixel_index2 >= 5681) && (pixel_index2 <= 5682)) || ((pixel_index2 >= 5684) && (pixel_index2 <= 5685)) || ((pixel_index2 >= 5690) && (pixel_index2 <= 5691)) || ((pixel_index2 >= 5693) && (pixel_index2 <= 5698)) || ((pixel_index2 >= 5700) && (pixel_index2 <= 5705)) || ((pixel_index2 >= 5707) && (pixel_index2 <= 5708)) || ((pixel_index2 >= 5710) && (pixel_index2 <= 5715)) || ((pixel_index2 >= 5721) && (pixel_index2 <= 5728)) || ((pixel_index2 >= 5730) && (pixel_index2 <= 5735)) || ((pixel_index2 >= 5737) && (pixel_index2 <= 5744)) || ((pixel_index2 >= 5746) && (pixel_index2 <= 5751)) || ((pixel_index2 >= 5769) && (pixel_index2 <= 5774)) || pixel_index2 == 5777 || pixel_index2 == 5781 || pixel_index2 == 5786 || ((pixel_index2 >= 5790) && (pixel_index2 <= 5793)) || ((pixel_index2 >= 5797) && (pixel_index2 <= 5800)) || pixel_index2 == 5803 || ((pixel_index2 >= 5807) && (pixel_index2 <= 5810)) || ((pixel_index2 >= 5818) && (pixel_index2 <= 5823)) || ((pixel_index2 >= 5827) && (pixel_index2 <= 5830)) || ((pixel_index2 >= 5834) && (pixel_index2 <= 5839)) || (pixel_index2 >= 5843) && (pixel_index2 <= 5846)) oled_data2 = 16'b1111010100010100;
                    else oled_data2 = 0;
                end
                1: begin
                    if (pixel_index2 == 97 || pixel_index2 == 99 || pixel_index2 == 101 || ((pixel_index2 >= 103) && (pixel_index2 <= 104)) || ((pixel_index2 >= 106) && (pixel_index2 <= 109)) || pixel_index2 == 111 || ((pixel_index2 >= 113) && (pixel_index2 <= 114)) || ((pixel_index2 >= 118) && (pixel_index2 <= 120)) || pixel_index2 == 195 || pixel_index2 == 197 || ((pixel_index2 >= 199) && (pixel_index2 <= 200)) || pixel_index2 == 202 || ((pixel_index2 >= 204) && (pixel_index2 <= 205)) || pixel_index2 == 207 || ((pixel_index2 >= 209) && (pixel_index2 <= 210)) || pixel_index2 == 213 || pixel_index2 == 289 || ((pixel_index2 >= 291) && (pixel_index2 <= 296)) || pixel_index2 == 298 || ((pixel_index2 >= 300) && (pixel_index2 <= 301)) || pixel_index2 == 303 || ((pixel_index2 >= 305) && (pixel_index2 <= 306)) || ((pixel_index2 >= 310) && (pixel_index2 <= 312)) || pixel_index2 == 385 || ((pixel_index2 >= 387) && (pixel_index2 <= 392)) || pixel_index2 == 394 || ((pixel_index2 >= 396) && (pixel_index2 <= 397)) || ((pixel_index2 >= 399) && (pixel_index2 <= 402)) || pixel_index2 == 408 || ((pixel_index2 >= 501) && (pixel_index2 <= 504)) || ((pixel_index2 >= 674) && (pixel_index2 <= 675)) || ((pixel_index2 >= 678) && (pixel_index2 <= 681)) || ((pixel_index2 >= 685) && (pixel_index2 <= 686)) || pixel_index2 == 688 || ((pixel_index2 >= 690) && (pixel_index2 <= 691)) || ((pixel_index2 >= 693) && (pixel_index2 <= 696)) || ((pixel_index2 >= 770) && (pixel_index2 <= 771)) || pixel_index2 == 774 || ((pixel_index2 >= 776) && (pixel_index2 <= 777)) || ((pixel_index2 >= 779) && (pixel_index2 <= 782)) || pixel_index2 == 784 || ((pixel_index2 >= 786) && (pixel_index2 <= 787)) || ((pixel_index2 >= 790) && (pixel_index2 <= 791)) || ((pixel_index2 >= 866) && (pixel_index2 <= 867)) || pixel_index2 == 870 || ((pixel_index2 >= 872) && (pixel_index2 <= 873)) || pixel_index2 == 875 || ((pixel_index2 >= 877) && (pixel_index2 <= 878)) || pixel_index2 == 880 || ((pixel_index2 >= 882) && (pixel_index2 <= 883)) || ((pixel_index2 >= 886) && (pixel_index2 <= 887)) || ((pixel_index2 >= 895) && (pixel_index2 <= 896)) || ((pixel_index2 >= 899) && (pixel_index2 <= 900)) || ((pixel_index2 >= 903) && (pixel_index2 <= 904)) || ((pixel_index2 >= 907) && (pixel_index2 <= 908)) || ((pixel_index2 >= 911) && (pixel_index2 <= 912)) || ((pixel_index2 >= 915) && (pixel_index2 <= 916)) || ((pixel_index2 >= 919) && (pixel_index2 <= 920)) || ((pixel_index2 >= 923) && (pixel_index2 <= 924)) || ((pixel_index2 >= 927) && (pixel_index2 <= 928)) || ((pixel_index2 >= 931) && (pixel_index2 <= 932)) || ((pixel_index2 >= 935) && (pixel_index2 <= 936)) || ((pixel_index2 >= 939) && (pixel_index2 <= 940)) || ((pixel_index2 >= 943) && (pixel_index2 <= 944)) || ((pixel_index2 >= 947) && (pixel_index2 <= 948)) || ((pixel_index2 >= 951) && (pixel_index2 <= 952)) || ((pixel_index2 >= 955) && (pixel_index2 <= 956)) || ((pixel_index2 >= 961) && (pixel_index2 <= 964)) || pixel_index2 == 966 || ((pixel_index2 >= 968) && (pixel_index2 <= 969)) || ((pixel_index2 >= 971) && (pixel_index2 <= 974)) || ((pixel_index2 >= 976) && (pixel_index2 <= 979)) || ((pixel_index2 >= 981) && (pixel_index2 <= 984)) || pixel_index2 == 1155 || ((pixel_index2 >= 1159) && (pixel_index2 <= 1161)) || pixel_index2 == 1163 || ((pixel_index2 >= 1165) && (pixel_index2 <= 1166)) || pixel_index2 == 1168 || ((pixel_index2 >= 1170) && (pixel_index2 <= 1171)) || pixel_index2 == 1173 || ((pixel_index2 >= 1175) && (pixel_index2 <= 1176)) || pixel_index2 == 1254 || ((pixel_index2 >= 1256) && (pixel_index2 <= 1257)) || pixel_index2 == 1259 || ((pixel_index2 >= 1261) && (pixel_index2 <= 1262)) || ((pixel_index2 >= 1264) && (pixel_index2 <= 1267)) || ((pixel_index2 >= 1270) && (pixel_index2 <= 1272)) || pixel_index2 == 1350 || ((pixel_index2 >= 1352) && (pixel_index2 <= 1353)) || pixel_index2 == 1355 || ((pixel_index2 >= 1357) && (pixel_index2 <= 1358)) || pixel_index2 == 1360 || ((pixel_index2 >= 1362) && (pixel_index2 <= 1363)) || pixel_index2 == 1365 || ((pixel_index2 >= 1367) && (pixel_index2 <= 1368)) || ((pixel_index2 >= 1447) && (pixel_index2 <= 1449)) || ((pixel_index2 >= 1451) && (pixel_index2 <= 1454)) || ((pixel_index2 >= 1456) && (pixel_index2 <= 1459)) || ((pixel_index2 >= 1461) && (pixel_index2 <= 1464)) || ((pixel_index2 >= 1637) && (pixel_index2 <= 1638)) || ((pixel_index2 >= 1641) && (pixel_index2 <= 1644)) || ((pixel_index2 >= 1646) && (pixel_index2 <= 1649)) || ((pixel_index2 >= 1652) && (pixel_index2 <= 1654)) || pixel_index2 == 1732 || pixel_index2 == 1735 || pixel_index2 == 1740 || pixel_index2 == 1745 || pixel_index2 == 1747 || pixel_index2 == 1831 || pixel_index2 == 1836 || ((pixel_index2 >= 1839) && (pixel_index2 <= 1841)) || ((pixel_index2 >= 1844) && (pixel_index2 <= 1845)) || pixel_index2 == 1924 || pixel_index2 == 1927 || pixel_index2 == 1932 || pixel_index2 == 1937 || pixel_index2 == 1942 || ((pixel_index2 >= 2021) && (pixel_index2 <= 2022)) || pixel_index2 == 2028 || ((pixel_index2 >= 2030) && (pixel_index2 <= 2033)) || ((pixel_index2 >= 2035) && (pixel_index2 <= 2037)) || pixel_index2 == 2213 || pixel_index2 == 2216 || ((pixel_index2 >= 2219) && (pixel_index2 <= 2221)) || pixel_index2 == 2223 || pixel_index2 == 2226 || ((pixel_index2 >= 2228) && (pixel_index2 <= 2230)) || pixel_index2 == 2310 || pixel_index2 == 2312 || pixel_index2 == 2314 || pixel_index2 == 2319 || pixel_index2 == 2322 || pixel_index2 == 2325 || ((pixel_index2 >= 2406) && (pixel_index2 <= 2408)) || ((pixel_index2 >= 2411) && (pixel_index2 <= 2412)) || ((pixel_index2 >= 2415) && (pixel_index2 <= 2416)) || pixel_index2 == 2418 || pixel_index2 == 2421 || pixel_index2 == 2501 || pixel_index2 == 2504 || pixel_index2 == 2509 || pixel_index2 == 2511 || ((pixel_index2 >= 2513) && (pixel_index2 <= 2514)) || pixel_index2 == 2517 || ((pixel_index2 >= 2598) && (pixel_index2 <= 2600)) || ((pixel_index2 >= 2602) && (pixel_index2 <= 2604)) || pixel_index2 == 2607 || pixel_index2 == 2610 || ((pixel_index2 >= 2612) && (pixel_index2 <= 2614)) || pixel_index2 == 2788 || pixel_index2 == 2791 || ((pixel_index2 >= 2794) && (pixel_index2 <= 2795)) || ((pixel_index2 >= 2799) && (pixel_index2 <= 2800)) || ((pixel_index2 >= 2804) && (pixel_index2 <= 2805)) || pixel_index2 == 2885 || pixel_index2 == 2887 || pixel_index2 == 2889 || pixel_index2 == 2892 || pixel_index2 == 2894 || pixel_index2 == 2897 || pixel_index2 == 2899 || pixel_index2 == 2902 || ((pixel_index2 >= 2982) && (pixel_index2 <= 2983)) || pixel_index2 == 2988 || pixel_index2 == 2990 || pixel_index2 == 2993 || pixel_index2 == 2998 || pixel_index2 == 3077 || pixel_index2 == 3079 || pixel_index2 == 3081 || pixel_index2 == 3084 || pixel_index2 == 3086 || pixel_index2 == 3089 || pixel_index2 == 3091 || pixel_index2 == 3094 || ((pixel_index2 >= 3133) && (pixel_index2 <= 3134)) || pixel_index2 == 3172 || pixel_index2 == 3175 || ((pixel_index2 >= 3178) && (pixel_index2 <= 3179)) || ((pixel_index2 >= 3183) && (pixel_index2 <= 3184)) || ((pixel_index2 >= 3188) && (pixel_index2 <= 3189)) || pixel_index2 == 3228 || pixel_index2 == 3327 || ((pixel_index2 >= 3364) && (pixel_index2 <= 3367)) || ((pixel_index2 >= 3370) && (pixel_index2 <= 3372)) || ((pixel_index2 >= 3375) && (pixel_index2 <= 3376)) || ((pixel_index2 >= 3380) && (pixel_index2 <= 3382)) || pixel_index2 == 3463 || pixel_index2 == 3465 || pixel_index2 == 3468 || pixel_index2 == 3470 || pixel_index2 == 3473 || pixel_index2 == 3475 || pixel_index2 == 3478 || pixel_index2 == 3559 || ((pixel_index2 >= 3562) && (pixel_index2 <= 3564)) || pixel_index2 == 3566 || pixel_index2 == 3569 || ((pixel_index2 >= 3572) && (pixel_index2 <= 3574)) || ((pixel_index2 >= 3630) && (pixel_index2 <= 3631)) || pixel_index2 == 3655 || pixel_index2 == 3657 || pixel_index2 == 3660 || pixel_index2 == 3662 || pixel_index2 == 3665 || pixel_index2 == 3667 || pixel_index2 == 3670 || pixel_index2 == 3751 || ((pixel_index2 >= 3754) && (pixel_index2 <= 3756)) || pixel_index2 == 3758 || pixel_index2 == 3761 || ((pixel_index2 >= 3764) && (pixel_index2 <= 3766)) || ((pixel_index2 >= 3938) && (pixel_index2 <= 3939)) || pixel_index2 == 3942 || pixel_index2 == 3945 || ((pixel_index2 >= 3947) && (pixel_index2 <= 3950)) || pixel_index2 == 3952 || ((pixel_index2 >= 3954) && (pixel_index2 <= 3955)) || ((pixel_index2 >= 3959) && (pixel_index2 <= 3962)) || ((pixel_index2 >= 3964) && (pixel_index2 <= 3967)) || ((pixel_index2 >= 3969) && (pixel_index2 <= 3972)) || ((pixel_index2 >= 3974) && (pixel_index2 <= 3977)) || pixel_index2 == 3979 || ((pixel_index2 >= 3981) && (pixel_index2 <= 3982)) || ((pixel_index2 >= 3984) && (pixel_index2 <= 3986)) || ((pixel_index2 >= 4008) && (pixel_index2 <= 4009)) || ((pixel_index2 >= 4012) && (pixel_index2 <= 4015)) || ((pixel_index2 >= 4017) && (pixel_index2 <= 4020)) || ((pixel_index2 >= 4022) && (pixel_index2 <= 4025)) || pixel_index2 == 4027 || ((pixel_index2 >= 4029) && (pixel_index2 <= 4030)) || ((pixel_index2 >= 4034) && (pixel_index2 <= 4035)) || ((pixel_index2 >= 4039) && (pixel_index2 <= 4040)) || ((pixel_index2 >= 4045) && (pixel_index2 <= 4046)) || pixel_index2 == 4048 || ((pixel_index2 >= 4050) && (pixel_index2 <= 4051)) || ((pixel_index2 >= 4057) && (pixel_index2 <= 4058)) || ((pixel_index2 >= 4060) && (pixel_index2 <= 4061)) || pixel_index2 == 4065 || ((pixel_index2 >= 4067) && (pixel_index2 <= 4068)) || pixel_index2 == 4070 || ((pixel_index2 >= 4072) && (pixel_index2 <= 4073)) || ((pixel_index2 >= 4075) && (pixel_index2 <= 4078)) || ((pixel_index2 >= 4082) && (pixel_index2 <= 4083)) || ((pixel_index2 >= 4104) && (pixel_index2 <= 4105)) || ((pixel_index2 >= 4110) && (pixel_index2 <= 4111)) || ((pixel_index2 >= 4113) && (pixel_index2 <= 4114)) || ((pixel_index2 >= 4120) && (pixel_index2 <= 4121)) || ((pixel_index2 >= 4124) && (pixel_index2 <= 4126)) || ((pixel_index2 >= 4130) && (pixel_index2 <= 4131)) || ((pixel_index2 >= 4135) && (pixel_index2 <= 4136)) || ((pixel_index2 >= 4139) && (pixel_index2 <= 4140)) || pixel_index2 == 4142 || pixel_index2 == 4144 || ((pixel_index2 >= 4146) && (pixel_index2 <= 4147)) || ((pixel_index2 >= 4151) && (pixel_index2 <= 4152)) || pixel_index2 == 4154 || ((pixel_index2 >= 4157) && (pixel_index2 <= 4159)) || pixel_index2 == 4161 || ((pixel_index2 >= 4163) && (pixel_index2 <= 4164)) || pixel_index2 == 4166 || ((pixel_index2 >= 4168) && (pixel_index2 <= 4169)) || pixel_index2 == 4171 || ((pixel_index2 >= 4173) && (pixel_index2 <= 4174)) || ((pixel_index2 >= 4178) && (pixel_index2 <= 4179)) || ((pixel_index2 >= 4200) && (pixel_index2 <= 4201)) || ((pixel_index2 >= 4204) && (pixel_index2 <= 4205)) || pixel_index2 == 4207 || ((pixel_index2 >= 4210) && (pixel_index2 <= 4212)) || ((pixel_index2 >= 4214) && (pixel_index2 <= 4215)) || pixel_index2 == 4217 || pixel_index2 == 4219 || ((pixel_index2 >= 4221) && (pixel_index2 <= 4222)) || ((pixel_index2 >= 4225) && (pixel_index2 <= 4228)) || pixel_index2 == 4230 || pixel_index2 == 4233 || ((pixel_index2 >= 4235) && (pixel_index2 <= 4238)) || ((pixel_index2 >= 4240) && (pixel_index2 <= 4243)) || ((pixel_index2 >= 4247) && (pixel_index2 <= 4250)) || ((pixel_index2 >= 4252) && (pixel_index2 <= 4254)) || ((pixel_index2 >= 4257) && (pixel_index2 <= 4260)) || ((pixel_index2 >= 4262) && (pixel_index2 <= 4265)) || pixel_index2 == 4267 || ((pixel_index2 >= 4269) && (pixel_index2 <= 4270)) || ((pixel_index2 >= 4272) && (pixel_index2 <= 4274)) || ((pixel_index2 >= 4295) && (pixel_index2 <= 4298)) || ((pixel_index2 >= 4300) && (pixel_index2 <= 4303)) || ((pixel_index2 >= 4305) && (pixel_index2 <= 4307)) || ((pixel_index2 >= 4310) && (pixel_index2 <= 4313)) || ((pixel_index2 >= 4315) && (pixel_index2 <= 4318)) || pixel_index2 == 4802 || pixel_index2 == 4893 || pixel_index2 == 5762 || pixel_index2 == 5853) oled_data2 = 16'b1111011110011110;
                    else if (((pixel_index2 >= 124) && (pixel_index2 <= 190)) || ((pixel_index2 >= 220) && (pixel_index2 <= 221)) || pixel_index2 == 225 || pixel_index2 == 229 || pixel_index2 == 233 || pixel_index2 == 237 || pixel_index2 == 241 || pixel_index2 == 245 || pixel_index2 == 249 || pixel_index2 == 253 || pixel_index2 == 257 || pixel_index2 == 261 || pixel_index2 == 265 || pixel_index2 == 269 || pixel_index2 == 273 || pixel_index2 == 277 || pixel_index2 == 281 || ((pixel_index2 >= 285) && (pixel_index2 <= 286)) || ((pixel_index2 >= 316) && (pixel_index2 <= 317)) || pixel_index2 == 321 || pixel_index2 == 325 || pixel_index2 == 329 || pixel_index2 == 333 || pixel_index2 == 337 || pixel_index2 == 341 || pixel_index2 == 345 || pixel_index2 == 349 || pixel_index2 == 353 || pixel_index2 == 357 || pixel_index2 == 361 || pixel_index2 == 365 || pixel_index2 == 369 || pixel_index2 == 373 || pixel_index2 == 377 || ((pixel_index2 >= 381) && (pixel_index2 <= 382)) || ((pixel_index2 >= 412) && (pixel_index2 <= 413)) || pixel_index2 == 417 || pixel_index2 == 421 || pixel_index2 == 425 || pixel_index2 == 429 || pixel_index2 == 433 || pixel_index2 == 437 || pixel_index2 == 441 || pixel_index2 == 445 || pixel_index2 == 449 || pixel_index2 == 453 || pixel_index2 == 457 || pixel_index2 == 461 || pixel_index2 == 465 || pixel_index2 == 469 || pixel_index2 == 473 || ((pixel_index2 >= 477) && (pixel_index2 <= 478)) || ((pixel_index2 >= 508) && (pixel_index2 <= 509)) || pixel_index2 == 513 || pixel_index2 == 517 || pixel_index2 == 521 || pixel_index2 == 525 || pixel_index2 == 529 || pixel_index2 == 533 || pixel_index2 == 537 || pixel_index2 == 541 || pixel_index2 == 545 || pixel_index2 == 549 || pixel_index2 == 553 || pixel_index2 == 557 || pixel_index2 == 561 || pixel_index2 == 565 || pixel_index2 == 569 || ((pixel_index2 >= 573) && (pixel_index2 <= 574)) || ((pixel_index2 >= 604) && (pixel_index2 <= 605)) || pixel_index2 == 609 || pixel_index2 == 613 || pixel_index2 == 617 || pixel_index2 == 621 || pixel_index2 == 625 || pixel_index2 == 629 || pixel_index2 == 633 || pixel_index2 == 637 || pixel_index2 == 641 || pixel_index2 == 645 || pixel_index2 == 649 || pixel_index2 == 653 || pixel_index2 == 657 || pixel_index2 == 661 || pixel_index2 == 665 || ((pixel_index2 >= 669) && (pixel_index2 <= 670)) || ((pixel_index2 >= 700) && (pixel_index2 <= 701)) || pixel_index2 == 705 || pixel_index2 == 709 || pixel_index2 == 713 || pixel_index2 == 717 || pixel_index2 == 721 || pixel_index2 == 725 || pixel_index2 == 729 || pixel_index2 == 733 || pixel_index2 == 737 || pixel_index2 == 741 || pixel_index2 == 745 || pixel_index2 == 749 || pixel_index2 == 753 || pixel_index2 == 757 || pixel_index2 == 761 || ((pixel_index2 >= 765) && (pixel_index2 <= 766)) || ((pixel_index2 >= 796) && (pixel_index2 <= 862)) || ((pixel_index2 >= 892) && (pixel_index2 <= 894)) || ((pixel_index2 >= 897) && (pixel_index2 <= 898)) || ((pixel_index2 >= 901) && (pixel_index2 <= 902)) || ((pixel_index2 >= 905) && (pixel_index2 <= 906)) || ((pixel_index2 >= 909) && (pixel_index2 <= 910)) || ((pixel_index2 >= 913) && (pixel_index2 <= 914)) || ((pixel_index2 >= 917) && (pixel_index2 <= 918)) || ((pixel_index2 >= 921) && (pixel_index2 <= 922)) || ((pixel_index2 >= 925) && (pixel_index2 <= 926)) || ((pixel_index2 >= 929) && (pixel_index2 <= 930)) || ((pixel_index2 >= 933) && (pixel_index2 <= 934)) || ((pixel_index2 >= 937) && (pixel_index2 <= 938)) || ((pixel_index2 >= 941) && (pixel_index2 <= 942)) || ((pixel_index2 >= 945) && (pixel_index2 <= 946)) || ((pixel_index2 >= 949) && (pixel_index2 <= 950)) || ((pixel_index2 >= 953) && (pixel_index2 <= 954)) || ((pixel_index2 >= 957) && (pixel_index2 <= 958)) || ((pixel_index2 >= 988) && (pixel_index2 <= 1054)) || ((pixel_index2 >= 1084) && (pixel_index2 <= 1085)) || ((pixel_index2 >= 1087) && (pixel_index2 <= 1089)) || ((pixel_index2 >= 1091) && (pixel_index2 <= 1093)) || ((pixel_index2 >= 1095) && (pixel_index2 <= 1097)) || ((pixel_index2 >= 1099) && (pixel_index2 <= 1101)) || ((pixel_index2 >= 1103) && (pixel_index2 <= 1105)) || ((pixel_index2 >= 1107) && (pixel_index2 <= 1109)) || ((pixel_index2 >= 1111) && (pixel_index2 <= 1113)) || ((pixel_index2 >= 1115) && (pixel_index2 <= 1117)) || ((pixel_index2 >= 1119) && (pixel_index2 <= 1121)) || ((pixel_index2 >= 1123) && (pixel_index2 <= 1125)) || ((pixel_index2 >= 1127) && (pixel_index2 <= 1129)) || ((pixel_index2 >= 1131) && (pixel_index2 <= 1133)) || ((pixel_index2 >= 1135) && (pixel_index2 <= 1137)) || ((pixel_index2 >= 1139) && (pixel_index2 <= 1141)) || ((pixel_index2 >= 1143) && (pixel_index2 <= 1145)) || ((pixel_index2 >= 1147) && (pixel_index2 <= 1150)) || ((pixel_index2 >= 1182) && (pixel_index2 <= 1219)) || ((pixel_index2 >= 1240) && (pixel_index2 <= 1244)) || ((pixel_index2 >= 1278) && (pixel_index2 <= 1280)) || ((pixel_index2 >= 1283) && (pixel_index2 <= 1286)) || ((pixel_index2 >= 1290) && (pixel_index2 <= 1291)) || ((pixel_index2 >= 1293) && (pixel_index2 <= 1294)) || ((pixel_index2 >= 1314) && (pixel_index2 <= 1315)) || ((pixel_index2 >= 1336) && (pixel_index2 <= 1340)) || ((pixel_index2 >= 1374) && (pixel_index2 <= 1376)) || ((pixel_index2 >= 1378) && (pixel_index2 <= 1382)) || ((pixel_index2 >= 1386) && (pixel_index2 <= 1390)) || ((pixel_index2 >= 1410) && (pixel_index2 <= 1411)) || ((pixel_index2 >= 1432) && (pixel_index2 <= 1436)) || ((pixel_index2 >= 1470) && (pixel_index2 <= 1478)) || ((pixel_index2 >= 1482) && (pixel_index2 <= 1486)) || ((pixel_index2 >= 1506) && (pixel_index2 <= 1507)) || ((pixel_index2 >= 1528) && (pixel_index2 <= 1532)) || ((pixel_index2 >= 1566) && (pixel_index2 <= 1603)) || ((pixel_index2 >= 1624) && (pixel_index2 <= 1628)) || ((pixel_index2 >= 1662) && (pixel_index2 <= 1666)) || pixel_index2 == 1670 || pixel_index2 == 1674 || ((pixel_index2 >= 1678) && (pixel_index2 <= 1696)) || ((pixel_index2 >= 1698) && (pixel_index2 <= 1699)) || ((pixel_index2 >= 1720) && (pixel_index2 <= 1724)) || ((pixel_index2 >= 1758) && (pixel_index2 <= 1762)) || pixel_index2 == 1766 || pixel_index2 == 1770 || ((pixel_index2 >= 1774) && (pixel_index2 <= 1775)) || ((pixel_index2 >= 1777) && (pixel_index2 <= 1789)) || pixel_index2 == 1792 || ((pixel_index2 >= 1794) && (pixel_index2 <= 1795)) || pixel_index2 == 1816 || ((pixel_index2 >= 1818) && (pixel_index2 <= 1820)) || ((pixel_index2 >= 1854) && (pixel_index2 <= 1858)) || pixel_index2 == 1862 || pixel_index2 == 1866 || pixel_index2 == 1870 || ((pixel_index2 >= 1872) && (pixel_index2 <= 1878)) || ((pixel_index2 >= 1882) && (pixel_index2 <= 1888)) || ((pixel_index2 >= 1892) && (pixel_index2 <= 1913)) || ((pixel_index2 >= 1915) && (pixel_index2 <= 1916)) || ((pixel_index2 >= 1948) && (pixel_index2 <= 1973)) || pixel_index2 == 1988 || pixel_index2 == 1991 || ((pixel_index2 >= 1993) && (pixel_index2 <= 1994)) || pixel_index2 == 1996 || ((pixel_index2 >= 2000) && (pixel_index2 <= 2001)) || pixel_index2 == 2008 || ((pixel_index2 >= 2011) && (pixel_index2 <= 2014)) || ((pixel_index2 >= 2044) && (pixel_index2 <= 2046)) || ((pixel_index2 >= 2048) && (pixel_index2 <= 2054)) || ((pixel_index2 >= 2058) && (pixel_index2 <= 2069)) || ((pixel_index2 >= 2084) && (pixel_index2 <= 2085)) || pixel_index2 == 2089 || ((pixel_index2 >= 2091) && (pixel_index2 <= 2093)) || ((pixel_index2 >= 2095) && (pixel_index2 <= 2096)) || ((pixel_index2 >= 2104) && (pixel_index2 <= 2105)) || ((pixel_index2 >= 2107) && (pixel_index2 <= 2110)) || pixel_index2 == 2140 || pixel_index2 == 2142 || ((pixel_index2 >= 2144) && (pixel_index2 <= 2150)) || pixel_index2 == 2154 || ((pixel_index2 >= 2157) && (pixel_index2 <= 2168)) || pixel_index2 == 2178 || ((pixel_index2 >= 2180) && (pixel_index2 <= 2184)) || pixel_index2 == 2188 || ((pixel_index2 >= 2190) && (pixel_index2 <= 2192)) || ((pixel_index2 >= 2195) && (pixel_index2 <= 2197)) || ((pixel_index2 >= 2200) && (pixel_index2 <= 2206)) || ((pixel_index2 >= 2236) && (pixel_index2 <= 2238)) || ((pixel_index2 >= 2245) && (pixel_index2 <= 2246)) || pixel_index2 == 2250 || ((pixel_index2 >= 2252) && (pixel_index2 <= 2264)) || ((pixel_index2 >= 2274) && (pixel_index2 <= 2288)) || ((pixel_index2 >= 2291) && (pixel_index2 <= 2293)) || ((pixel_index2 >= 2296) && (pixel_index2 <= 2302)) || ((pixel_index2 >= 2332) && (pixel_index2 <= 2334)) || ((pixel_index2 >= 2341) && (pixel_index2 <= 2355)) || ((pixel_index2 >= 2374) && (pixel_index2 <= 2384)) || ((pixel_index2 >= 2392) && (pixel_index2 <= 2398)) || ((pixel_index2 >= 2428) && (pixel_index2 <= 2437)) || ((pixel_index2 >= 2443) && (pixel_index2 <= 2451)) || ((pixel_index2 >= 2470) && (pixel_index2 <= 2480)) || ((pixel_index2 >= 2487) && (pixel_index2 <= 2494)) || ((pixel_index2 >= 2526) && (pixel_index2 <= 2532)) || ((pixel_index2 >= 2540) && (pixel_index2 <= 2547)) || pixel_index2 == 2566 || ((pixel_index2 >= 2580) && (pixel_index2 <= 2588)) || ((pixel_index2 >= 2622) && (pixel_index2 <= 2626)) || pixel_index2 == 2636 || ((pixel_index2 >= 2639) && (pixel_index2 <= 2644)) || ((pixel_index2 >= 2647) && (pixel_index2 <= 2648)) || pixel_index2 == 2659 || ((pixel_index2 >= 2661) && (pixel_index2 <= 2662)) || ((pixel_index2 >= 2676) && (pixel_index2 <= 2684)) || ((pixel_index2 >= 2718) && (pixel_index2 <= 2721)) || pixel_index2 == 2732 || ((pixel_index2 >= 2735) && (pixel_index2 <= 2742)) || ((pixel_index2 >= 2756) && (pixel_index2 <= 2758)) || ((pixel_index2 >= 2772) && (pixel_index2 <= 2780)) || ((pixel_index2 >= 2814) && (pixel_index2 <= 2817)) || pixel_index2 == 2828 || ((pixel_index2 >= 2831) && (pixel_index2 <= 2838)) || ((pixel_index2 >= 2842) && (pixel_index2 <= 2848)) || ((pixel_index2 >= 2852) && (pixel_index2 <= 2859)) || ((pixel_index2 >= 2866) && (pixel_index2 <= 2876)) || ((pixel_index2 >= 2910) && (pixel_index2 <= 2913)) || pixel_index2 == 2924 || ((pixel_index2 >= 2927) && (pixel_index2 <= 2935)) || ((pixel_index2 >= 2938) && (pixel_index2 <= 2944)) || ((pixel_index2 >= 2947) && (pixel_index2 <= 2955)) || pixel_index2 == 2962 || ((pixel_index2 >= 2964) && (pixel_index2 <= 2972)) || ((pixel_index2 >= 3006) && (pixel_index2 <= 3013)) || ((pixel_index2 >= 3019) && (pixel_index2 <= 3021)) || ((pixel_index2 >= 3023) && (pixel_index2 <= 3032)) || ((pixel_index2 >= 3042) && (pixel_index2 <= 3051)) || ((pixel_index2 >= 3058) && (pixel_index2 <= 3060)) || pixel_index2 == 3063 || ((pixel_index2 >= 3065) && (pixel_index2 <= 3068)) || ((pixel_index2 >= 3102) && (pixel_index2 <= 3104)) || pixel_index2 == 3107 || ((pixel_index2 >= 3117) && (pixel_index2 <= 3123)) || ((pixel_index2 >= 3143) && (pixel_index2 <= 3147)) || ((pixel_index2 >= 3154) && (pixel_index2 <= 3155)) || pixel_index2 == 3159 || ((pixel_index2 >= 3161) && (pixel_index2 <= 3164)) || ((pixel_index2 >= 3198) && (pixel_index2 <= 3200)) || ((pixel_index2 >= 3202) && (pixel_index2 <= 3203)) || ((pixel_index2 >= 3213) && (pixel_index2 <= 3216)) || ((pixel_index2 >= 3218) && (pixel_index2 <= 3219)) || ((pixel_index2 >= 3239) && (pixel_index2 <= 3243)) || ((pixel_index2 >= 3250) && (pixel_index2 <= 3251)) || ((pixel_index2 >= 3255) && (pixel_index2 <= 3260)) || ((pixel_index2 >= 3292) && (pixel_index2 <= 3299)) || ((pixel_index2 >= 3309) && (pixel_index2 <= 3312)) || ((pixel_index2 >= 3314) && (pixel_index2 <= 3315)) || ((pixel_index2 >= 3335) && (pixel_index2 <= 3337)) || pixel_index2 == 3339 || ((pixel_index2 >= 3346) && (pixel_index2 <= 3347)) || ((pixel_index2 >= 3351) && (pixel_index2 <= 3352)) || ((pixel_index2 >= 3354) && (pixel_index2 <= 3358)) || ((pixel_index2 >= 3388) && (pixel_index2 <= 3393)) || pixel_index2 == 3395 || ((pixel_index2 >= 3405) && (pixel_index2 <= 3407)) || ((pixel_index2 >= 3409) && (pixel_index2 <= 3411)) || ((pixel_index2 >= 3431) && (pixel_index2 <= 3432)) || ((pixel_index2 >= 3434) && (pixel_index2 <= 3435)) || ((pixel_index2 >= 3438) && (pixel_index2 <= 3443)) || ((pixel_index2 >= 3447) && (pixel_index2 <= 3448)) || ((pixel_index2 >= 3450) && (pixel_index2 <= 3454)) || ((pixel_index2 >= 3484) && (pixel_index2 <= 3487)) || pixel_index2 == 3489 || pixel_index2 == 3491 || ((pixel_index2 >= 3501) && (pixel_index2 <= 3502)) || ((pixel_index2 >= 3505) && (pixel_index2 <= 3507)) || ((pixel_index2 >= 3527) && (pixel_index2 <= 3531)) || ((pixel_index2 >= 3538) && (pixel_index2 <= 3539)) || ((pixel_index2 >= 3543) && (pixel_index2 <= 3544)) || ((pixel_index2 >= 3546) && (pixel_index2 <= 3550)) || ((pixel_index2 >= 3580) && (pixel_index2 <= 3587)) || ((pixel_index2 >= 3597) && (pixel_index2 <= 3603)) || ((pixel_index2 >= 3623) && (pixel_index2 <= 3628)) || ((pixel_index2 >= 3633) && (pixel_index2 <= 3635)) || ((pixel_index2 >= 3639) && (pixel_index2 <= 3646)) || ((pixel_index2 >= 4620) && (pixel_index2 <= 4692)) || ((pixel_index2 >= 4707) && (pixel_index2 <= 4796)) || ((pixel_index2 >= 4803) && (pixel_index2 <= 4812)) || ((pixel_index2 >= 4814) && (pixel_index2 <= 4817)) || ((pixel_index2 >= 4819) && (pixel_index2 <= 4820)) || ((pixel_index2 >= 4827) && (pixel_index2 <= 4829)) || ((pixel_index2 >= 4834) && (pixel_index2 <= 4835)) || ((pixel_index2 >= 4838) && (pixel_index2 <= 4839)) || ((pixel_index2 >= 4841) && (pixel_index2 <= 4843)) || ((pixel_index2 >= 4845) && (pixel_index2 <= 4846)) || ((pixel_index2 >= 4851) && (pixel_index2 <= 4861)) || ((pixel_index2 >= 4863) && (pixel_index2 <= 4865)) || ((pixel_index2 >= 4868) && (pixel_index2 <= 4869)) || ((pixel_index2 >= 4871) && (pixel_index2 <= 4873)) || ((pixel_index2 >= 4880) && (pixel_index2 <= 4882)) || ((pixel_index2 >= 4887) && (pixel_index2 <= 4892)) || ((pixel_index2 >= 4899) && (pixel_index2 <= 4907)) || ((pixel_index2 >= 4910) && (pixel_index2 <= 4912)) || pixel_index2 == 4915 || pixel_index2 == 4924 || pixel_index2 == 4931 || pixel_index2 == 4935 || pixel_index2 == 4938 || pixel_index2 == 4941 || ((pixel_index2 >= 4948) && (pixel_index2 <= 4956)) || ((pixel_index2 >= 4959) && (pixel_index2 <= 4961)) || pixel_index2 == 4965 || pixel_index2 == 4968 || pixel_index2 == 4977 || ((pixel_index2 >= 4984) && (pixel_index2 <= 4988)) || ((pixel_index2 >= 4994) && (pixel_index2 <= 5003)) || ((pixel_index2 >= 5006) && (pixel_index2 <= 5008)) || pixel_index2 == 5011 || pixel_index2 == 5020 || pixel_index2 == 5027 || pixel_index2 == 5034 || pixel_index2 == 5037 || ((pixel_index2 >= 5044) && (pixel_index2 <= 5052)) || ((pixel_index2 >= 5055) && (pixel_index2 <= 5057)) || pixel_index2 == 5064 || pixel_index2 == 5073 || ((pixel_index2 >= 5080) && (pixel_index2 <= 5085)) || ((pixel_index2 >= 5090) && (pixel_index2 <= 5099)) || ((pixel_index2 >= 5102) && (pixel_index2 <= 5104)) || pixel_index2 == 5107 || ((pixel_index2 >= 5111) && (pixel_index2 <= 5112)) || ((pixel_index2 >= 5116) && (pixel_index2 <= 5119)) || ((pixel_index2 >= 5123) && (pixel_index2 <= 5124)) || pixel_index2 == 5130 || ((pixel_index2 >= 5133) && (pixel_index2 <= 5136)) || ((pixel_index2 >= 5140) && (pixel_index2 <= 5148)) || ((pixel_index2 >= 5151) && (pixel_index2 <= 5154)) || pixel_index2 == 5160 || ((pixel_index2 >= 5164) && (pixel_index2 <= 5165)) || pixel_index2 == 5169 || ((pixel_index2 >= 5173) && (pixel_index2 <= 5181)) || ((pixel_index2 >= 5186) && (pixel_index2 <= 5195)) || ((pixel_index2 >= 5198) && (pixel_index2 <= 5200)) || pixel_index2 == 5203 || ((pixel_index2 >= 5206) && (pixel_index2 <= 5209)) || ((pixel_index2 >= 5212) && (pixel_index2 <= 5216)) || ((pixel_index2 >= 5219) && (pixel_index2 <= 5220)) || pixel_index2 == 5226 || ((pixel_index2 >= 5229) && (pixel_index2 <= 5233)) || ((pixel_index2 >= 5236) && (pixel_index2 <= 5244)) || ((pixel_index2 >= 5247) && (pixel_index2 <= 5250)) || pixel_index2 == 5256 || ((pixel_index2 >= 5259) && (pixel_index2 <= 5262)) || pixel_index2 == 5265 || ((pixel_index2 >= 5271) && (pixel_index2 <= 5277)) || ((pixel_index2 >= 5282) && (pixel_index2 <= 5291)) || ((pixel_index2 >= 5294) && (pixel_index2 <= 5296)) || pixel_index2 == 5299 || ((pixel_index2 >= 5302) && (pixel_index2 <= 5305)) || ((pixel_index2 >= 5308) && (pixel_index2 <= 5312)) || pixel_index2 == 5315 || pixel_index2 == 5322 || ((pixel_index2 >= 5325) && (pixel_index2 <= 5329)) || ((pixel_index2 >= 5332) && (pixel_index2 <= 5340)) || ((pixel_index2 >= 5343) && (pixel_index2 <= 5345)) || pixel_index2 == 5352 || ((pixel_index2 >= 5355) && (pixel_index2 <= 5358)) || pixel_index2 == 5361 || ((pixel_index2 >= 5368) && (pixel_index2 <= 5373)) || ((pixel_index2 >= 5378) && (pixel_index2 <= 5387)) || ((pixel_index2 >= 5390) && (pixel_index2 <= 5392)) || pixel_index2 == 5395 || ((pixel_index2 >= 5398) && (pixel_index2 <= 5401)) || ((pixel_index2 >= 5404) && (pixel_index2 <= 5408)) || pixel_index2 == 5411 || pixel_index2 == 5415 || pixel_index2 == 5418 || ((pixel_index2 >= 5421) && (pixel_index2 <= 5425)) || ((pixel_index2 >= 5428) && (pixel_index2 <= 5436)) || ((pixel_index2 >= 5439) && (pixel_index2 <= 5441)) || pixel_index2 == 5445 || pixel_index2 == 5448 || ((pixel_index2 >= 5451) && (pixel_index2 <= 5454)) || ((pixel_index2 >= 5457) && (pixel_index2 <= 5458)) || ((pixel_index2 >= 5464) && (pixel_index2 <= 5469)) || ((pixel_index2 >= 5474) && (pixel_index2 <= 5483)) || ((pixel_index2 >= 5486) && (pixel_index2 <= 5488)) || pixel_index2 == 5491 || ((pixel_index2 >= 5494) && (pixel_index2 <= 5497)) || ((pixel_index2 >= 5500) && (pixel_index2 <= 5503)) || pixel_index2 == 5507 || ((pixel_index2 >= 5510) && (pixel_index2 <= 5511)) || pixel_index2 == 5514 || ((pixel_index2 >= 5517) && (pixel_index2 <= 5520)) || ((pixel_index2 >= 5524) && (pixel_index2 <= 5532)) || ((pixel_index2 >= 5535) && (pixel_index2 <= 5537)) || ((pixel_index2 >= 5540) && (pixel_index2 <= 5541)) || pixel_index2 == 5544 || ((pixel_index2 >= 5548) && (pixel_index2 <= 5549)) || ((pixel_index2 >= 5553) && (pixel_index2 <= 5556)) || ((pixel_index2 >= 5560) && (pixel_index2 <= 5565)) || ((pixel_index2 >= 5570) && (pixel_index2 <= 5575)) || pixel_index2 == 5584 || pixel_index2 == 5587 || ((pixel_index2 >= 5590) && (pixel_index2 <= 5593)) || pixel_index2 == 5596 || pixel_index2 == 5603 || pixel_index2 == 5610 || pixel_index2 == 5613 || ((pixel_index2 >= 5620) && (pixel_index2 <= 5624)) || pixel_index2 == 5633 || pixel_index2 == 5640 || pixel_index2 == 5649 || ((pixel_index2 >= 5656) && (pixel_index2 <= 5661)) || ((pixel_index2 >= 5667) && (pixel_index2 <= 5671)) || pixel_index2 == 5680 || pixel_index2 == 5683 || ((pixel_index2 >= 5686) && (pixel_index2 <= 5689)) || pixel_index2 == 5692 || pixel_index2 == 5699 || pixel_index2 == 5706 || pixel_index2 == 5709 || ((pixel_index2 >= 5716) && (pixel_index2 <= 5720)) || pixel_index2 == 5729 || pixel_index2 == 5736 || pixel_index2 == 5745 || ((pixel_index2 >= 5752) && (pixel_index2 <= 5756)) || ((pixel_index2 >= 5763) && (pixel_index2 <= 5768)) || ((pixel_index2 >= 5775) && (pixel_index2 <= 5776)) || ((pixel_index2 >= 5778) && (pixel_index2 <= 5780)) || ((pixel_index2 >= 5782) && (pixel_index2 <= 5785)) || ((pixel_index2 >= 5787) && (pixel_index2 <= 5789)) || ((pixel_index2 >= 5794) && (pixel_index2 <= 5796)) || ((pixel_index2 >= 5801) && (pixel_index2 <= 5802)) || ((pixel_index2 >= 5804) && (pixel_index2 <= 5806)) || ((pixel_index2 >= 5811) && (pixel_index2 <= 5817)) || ((pixel_index2 >= 5824) && (pixel_index2 <= 5826)) || ((pixel_index2 >= 5831) && (pixel_index2 <= 5833)) || ((pixel_index2 >= 5840) && (pixel_index2 <= 5842)) || ((pixel_index2 >= 5847) && (pixel_index2 <= 5852)) || (pixel_index2 >= 5868) && (pixel_index2 <= 5940)) oled_data2 = 16'b0000000000001010;
                    else if (pixel_index2 == 511 || pixel_index2 == 515 || pixel_index2 == 519 || pixel_index2 == 523 || pixel_index2 == 527 || pixel_index2 == 531 || pixel_index2 == 535 || pixel_index2 == 539 || pixel_index2 == 543 || pixel_index2 == 547 || pixel_index2 == 551 || pixel_index2 == 555 || pixel_index2 == 559 || pixel_index2 == 563 || pixel_index2 == 567 || pixel_index2 == 571 || pixel_index2 == 607 || pixel_index2 == 611 || pixel_index2 == 615 || pixel_index2 == 619 || pixel_index2 == 623 || pixel_index2 == 627 || pixel_index2 == 631 || pixel_index2 == 635 || pixel_index2 == 639 || pixel_index2 == 643 || pixel_index2 == 647 || pixel_index2 == 651 || pixel_index2 == 655 || pixel_index2 == 659 || pixel_index2 == 663 || pixel_index2 == 667 || pixel_index2 == 3488) oled_data2 = 16'b1010000000000000;
                    else if (pixel_index2 == 1086 || pixel_index2 == 1114 || pixel_index2 == 1118 || pixel_index2 == 1122 || pixel_index2 == 1126 || pixel_index2 == 1130 || pixel_index2 == 1134 || pixel_index2 == 1138 || pixel_index2 == 1142 || pixel_index2 == 1146) oled_data2 = 16'b0000001010000000;
                    else if (pixel_index2 == 1090 || pixel_index2 == 1094 || pixel_index2 == 1098 || pixel_index2 == 1102 || pixel_index2 == 1106 || pixel_index2 == 1110 || pixel_index2 == 1287 || pixel_index2 == 1289 || pixel_index2 == 1479 || pixel_index2 == 1481 || pixel_index2 == 1667 || pixel_index2 == 1669 || pixel_index2 == 1671 || pixel_index2 == 1673 || pixel_index2 == 1675 || pixel_index2 == 1677 || pixel_index2 == 1859 || pixel_index2 == 1861 || pixel_index2 == 1863 || pixel_index2 == 1865 || pixel_index2 == 1867 || pixel_index2 == 1869 || ((pixel_index2 >= 1879) && (pixel_index2 <= 1881)) || ((pixel_index2 >= 1889) && (pixel_index2 <= 1891)) || ((pixel_index2 >= 1975) && (pixel_index2 <= 1987)) || ((pixel_index2 >= 2002) && (pixel_index2 <= 2007)) || pixel_index2 == 2055 || pixel_index2 == 2057 || ((pixel_index2 >= 2072) && (pixel_index2 <= 2073)) || ((pixel_index2 >= 2081) && (pixel_index2 <= 2082)) || ((pixel_index2 >= 2097) && (pixel_index2 <= 2103)) || pixel_index2 == 2169 || pixel_index2 == 2177 || ((pixel_index2 >= 2193) && (pixel_index2 <= 2194)) || ((pixel_index2 >= 2198) && (pixel_index2 <= 2199)) || pixel_index2 == 2239 || ((pixel_index2 >= 2241) && (pixel_index2 <= 2242)) || pixel_index2 == 2244 || pixel_index2 == 2247 || pixel_index2 == 2249 || pixel_index2 == 2265 || pixel_index2 == 2273 || ((pixel_index2 >= 2289) && (pixel_index2 <= 2290)) || ((pixel_index2 >= 2294) && (pixel_index2 <= 2295)) || pixel_index2 == 2335 || pixel_index2 == 2337 || pixel_index2 == 2339 || ((pixel_index2 >= 2356) && (pixel_index2 <= 2361)) || ((pixel_index2 >= 2369) && (pixel_index2 <= 2373)) || ((pixel_index2 >= 2385) && (pixel_index2 <= 2391)) || ((pixel_index2 >= 2438) && (pixel_index2 <= 2442)) || ((pixel_index2 >= 2452) && (pixel_index2 <= 2457)) || ((pixel_index2 >= 2465) && (pixel_index2 <= 2469)) || ((pixel_index2 >= 2481) && (pixel_index2 <= 2486)) || pixel_index2 == 2533 || pixel_index2 == 2539 || pixel_index2 == 2549 || ((pixel_index2 >= 2552) && (pixel_index2 <= 2553)) || pixel_index2 == 2561 || ((pixel_index2 >= 2564) && (pixel_index2 <= 2565)) || ((pixel_index2 >= 2627) && (pixel_index2 <= 2629)) || pixel_index2 == 2635 || ((pixel_index2 >= 2637) && (pixel_index2 <= 2638)) || pixel_index2 == 2649 || pixel_index2 == 2657 || ((pixel_index2 >= 2722) && (pixel_index2 <= 2725)) || pixel_index2 == 2731 || ((pixel_index2 >= 2733) && (pixel_index2 <= 2734)) || ((pixel_index2 >= 2743) && (pixel_index2 <= 2755)) || ((pixel_index2 >= 2818) && (pixel_index2 <= 2821)) || pixel_index2 == 2827 || ((pixel_index2 >= 2829) && (pixel_index2 <= 2830)) || ((pixel_index2 >= 2839) && (pixel_index2 <= 2841)) || ((pixel_index2 >= 2849) && (pixel_index2 <= 2851)) || ((pixel_index2 >= 2914) && (pixel_index2 <= 2917)) || pixel_index2 == 2923 || pixel_index2 == 2936 || pixel_index2 == 2945 || pixel_index2 == 2963 || ((pixel_index2 >= 3014) && (pixel_index2 <= 3018)) || ((pixel_index2 >= 3061) && (pixel_index2 <= 3062)) || pixel_index2 == 3064 || ((pixel_index2 >= 3108) && (pixel_index2 <= 3116)) || pixel_index2 == 3160 || ((pixel_index2 >= 3204) && (pixel_index2 <= 3212)) || ((pixel_index2 >= 3300) && (pixel_index2 <= 3308)) || pixel_index2 == 3317 || ((pixel_index2 >= 3319) && (pixel_index2 <= 3320)) || ((pixel_index2 >= 3330) && (pixel_index2 <= 3331)) || pixel_index2 == 3333 || pixel_index2 == 3338 || ((pixel_index2 >= 3396) && (pixel_index2 <= 3404)) || pixel_index2 == 3433 || ((pixel_index2 >= 3436) && (pixel_index2 <= 3437)) || ((pixel_index2 >= 3492) && (pixel_index2 <= 3500)) || ((pixel_index2 >= 3588) && (pixel_index2 <= 3596)) || ((pixel_index2 >= 3684) && (pixel_index2 <= 3692)) || ((pixel_index2 >= 3724) && (pixel_index2 <= 3729)) || ((pixel_index2 >= 3820) && (pixel_index2 <= 3825)) || ((pixel_index2 >= 3893) && (pixel_index2 <= 3894)) || ((pixel_index2 >= 3897) && (pixel_index2 <= 3905)) || ((pixel_index2 >= 3908) && (pixel_index2 <= 3909)) || ((pixel_index2 >= 3989) && (pixel_index2 <= 3990)) || ((pixel_index2 >= 3994) && (pixel_index2 <= 4000)) || ((pixel_index2 >= 4004) && (pixel_index2 <= 4005)) || ((pixel_index2 >= 4085) && (pixel_index2 <= 4086)) || ((pixel_index2 >= 4090) && (pixel_index2 <= 4096)) || ((pixel_index2 >= 4100) && (pixel_index2 <= 4101)) || pixel_index2 == 4706 || pixel_index2 == 4797 || pixel_index2 == 5666 || pixel_index2 == 5757) oled_data2 = 16'b0101001010001010;
                    else if (((pixel_index2 >= 1281) && (pixel_index2 <= 1282)) || pixel_index2 == 1292 || pixel_index2 == 1295 || ((pixel_index2 >= 1297) && (pixel_index2 <= 1299)) || pixel_index2 == 1302 || ((pixel_index2 >= 1304) && (pixel_index2 <= 1305)) || pixel_index2 == 1307 || pixel_index2 == 1309 || pixel_index2 == 1311 || pixel_index2 == 1313 || pixel_index2 == 1377 || ((pixel_index2 >= 1392) && (pixel_index2 <= 1395)) || ((pixel_index2 >= 1397) && (pixel_index2 <= 1399)) || pixel_index2 == 1401 || ((pixel_index2 >= 1403) && (pixel_index2 <= 1404)) || pixel_index2 == 1406 || pixel_index2 == 1409 || ((pixel_index2 >= 1487) && (pixel_index2 <= 1488)) || pixel_index2 == 1490 || pixel_index2 == 1493 || pixel_index2 == 1495 || pixel_index2 == 1497 || ((pixel_index2 >= 1499) && (pixel_index2 <= 1500)) || ((pixel_index2 >= 1502) && (pixel_index2 <= 1503)) || pixel_index2 == 1505 || pixel_index2 == 1697 || pixel_index2 == 1776 || ((pixel_index2 >= 1790) && (pixel_index2 <= 1791)) || pixel_index2 == 1793 || pixel_index2 == 1817 || pixel_index2 == 1871 || pixel_index2 == 1914 || pixel_index2 == 1974 || ((pixel_index2 >= 1989) && (pixel_index2 <= 1990)) || pixel_index2 == 1992 || pixel_index2 == 1995 || ((pixel_index2 >= 1997) && (pixel_index2 <= 1999)) || ((pixel_index2 >= 2009) && (pixel_index2 <= 2010)) || pixel_index2 == 2047 || ((pixel_index2 >= 2070) && (pixel_index2 <= 2071)) || pixel_index2 == 2083 || ((pixel_index2 >= 2086) && (pixel_index2 <= 2088)) || pixel_index2 == 2090 || pixel_index2 == 2094 || pixel_index2 == 2106 || pixel_index2 == 2141 || pixel_index2 == 2143 || ((pixel_index2 >= 2155) && (pixel_index2 <= 2156)) || pixel_index2 == 2179 || ((pixel_index2 >= 2185) && (pixel_index2 <= 2187)) || pixel_index2 == 2189 || pixel_index2 == 2240 || pixel_index2 == 2243 || pixel_index2 == 2251 || pixel_index2 == 2336 || pixel_index2 == 2338 || pixel_index2 == 2340 || pixel_index2 == 2548 || ((pixel_index2 >= 2550) && (pixel_index2 <= 2551)) || ((pixel_index2 >= 2562) && (pixel_index2 <= 2563)) || ((pixel_index2 >= 2567) && (pixel_index2 <= 2579)) || ((pixel_index2 >= 2645) && (pixel_index2 <= 2646)) || pixel_index2 == 2658 || pixel_index2 == 2660 || ((pixel_index2 >= 2663) && (pixel_index2 <= 2675)) || ((pixel_index2 >= 2759) && (pixel_index2 <= 2771)) || ((pixel_index2 >= 2925) && (pixel_index2 <= 2926)) || pixel_index2 == 2937 || pixel_index2 == 2946 || pixel_index2 == 3022 || ((pixel_index2 >= 3105) && (pixel_index2 <= 3106)) || pixel_index2 == 3201 || pixel_index2 == 3217 || ((pixel_index2 >= 3230) && (pixel_index2 <= 3231)) || pixel_index2 == 3313 || pixel_index2 == 3324 || pixel_index2 == 3408 || ((pixel_index2 >= 3421) && (pixel_index2 <= 3422)) || ((pixel_index2 >= 3503) && (pixel_index2 <= 3504)) || ((pixel_index2 >= 3533) && (pixel_index2 <= 3536)) || pixel_index2 == 3629 || pixel_index2 == 3632) oled_data2 = 16'b1010010100010100;
                    else if (pixel_index2 == 1296 || ((pixel_index2 >= 1300) && (pixel_index2 <= 1301)) || pixel_index2 == 1303 || pixel_index2 == 1306 || pixel_index2 == 1308 || pixel_index2 == 1310 || pixel_index2 == 1312 || pixel_index2 == 1391 || pixel_index2 == 1396 || pixel_index2 == 1400 || pixel_index2 == 1402 || pixel_index2 == 1405 || ((pixel_index2 >= 1407) && (pixel_index2 <= 1408)) || pixel_index2 == 1489 || ((pixel_index2 >= 1491) && (pixel_index2 <= 1492)) || pixel_index2 == 1494 || pixel_index2 == 1496 || pixel_index2 == 1498 || pixel_index2 == 1501 || pixel_index2 == 1504 || pixel_index2 == 3353 || pixel_index2 == 3449 || pixel_index2 == 3545) oled_data2 = 16'b0101001010010100;
                    else if (((pixel_index2 >= 1317) && (pixel_index2 <= 1319)) || pixel_index2 == 1324 || ((pixel_index2 >= 1327) && (pixel_index2 <= 1329)) || ((pixel_index2 >= 1332) && (pixel_index2 <= 1334)) || pixel_index2 == 1415 || pixel_index2 == 1420 || pixel_index2 == 1425 || pixel_index2 == 1428 || ((pixel_index2 >= 1509) && (pixel_index2 <= 1511)) || ((pixel_index2 >= 1514) && (pixel_index2 <= 1516)) || ((pixel_index2 >= 1519) && (pixel_index2 <= 1521)) || ((pixel_index2 >= 1524) && (pixel_index2 <= 1526)) || pixel_index2 == 1607 || pixel_index2 == 1617 || pixel_index2 == 1622 || pixel_index2 == 1703 || pixel_index2 == 1713 || (pixel_index2 >= 1716) && (pixel_index2 <= 1718)) oled_data2 = 16'b1010000000001010;
                    else if (pixel_index2 == 3229 || (pixel_index2 >= 3325) && (pixel_index2 <= 3326)) oled_data2 = 16'b0101010100001010;
                    else if (pixel_index2 == 3253 || pixel_index2 == 3349) oled_data2 = 16'b0000010100000000;
                    else if (pixel_index2 == 3394 || pixel_index2 == 3490) oled_data2 = 16'b0000000000010100;
                    else if (pixel_index2 == 3532 || pixel_index2 == 3537) oled_data2 = 16'b0101000000000000;
                    else if (((pixel_index2 >= 4423) && (pixel_index2 <= 4505)) || ((pixel_index2 >= 4513) && (pixel_index2 <= 4518)) || (pixel_index2 >= 4602) && (pixel_index2 <= 4606)) oled_data2 = 16'b0000001010011110;
                    else if (((pixel_index2 >= 4519) && (pixel_index2 <= 4601)) || ((pixel_index2 >= 4609) && (pixel_index2 <= 4619)) || ((pixel_index2 >= 4693) && (pixel_index2 <= 4702)) || pixel_index2 == 4705 || pixel_index2 == 4798 || pixel_index2 == 4801 || pixel_index2 == 4894 || ((pixel_index2 >= 4897) && (pixel_index2 <= 4898)) || ((pixel_index2 >= 4989) && (pixel_index2 <= 4990)) || pixel_index2 == 4993 || pixel_index2 == 5086 || pixel_index2 == 5089 || pixel_index2 == 5182 || pixel_index2 == 5185 || pixel_index2 == 5278 || pixel_index2 == 5281 || pixel_index2 == 5374 || pixel_index2 == 5377 || pixel_index2 == 5470 || pixel_index2 == 5473 || pixel_index2 == 5566 || pixel_index2 == 5569 || pixel_index2 == 5662 || pixel_index2 == 5665 || pixel_index2 == 5758 || pixel_index2 == 5761 || pixel_index2 == 5854 || ((pixel_index2 >= 5857) && (pixel_index2 <= 5867)) || ((pixel_index2 >= 5941) && (pixel_index2 <= 5950)) || (pixel_index2 >= 5959) && (pixel_index2 <= 6041)) oled_data2 = 16'b0000001010010100;
                    else if (pixel_index2 == 4813 || pixel_index2 == 4818 || ((pixel_index2 >= 4821) && (pixel_index2 <= 4826)) || ((pixel_index2 >= 4830) && (pixel_index2 <= 4833)) || ((pixel_index2 >= 4836) && (pixel_index2 <= 4837)) || pixel_index2 == 4840 || pixel_index2 == 4844 || ((pixel_index2 >= 4847) && (pixel_index2 <= 4850)) || pixel_index2 == 4862 || ((pixel_index2 >= 4866) && (pixel_index2 <= 4867)) || pixel_index2 == 4870 || ((pixel_index2 >= 4874) && (pixel_index2 <= 4879)) || ((pixel_index2 >= 4883) && (pixel_index2 <= 4886)) || pixel_index2 == 4908 || pixel_index2 == 4913 || pixel_index2 == 4916 || pixel_index2 == 4923 || pixel_index2 == 4925 || pixel_index2 == 4930 || pixel_index2 == 4934 || pixel_index2 == 4937 || pixel_index2 == 4939 || pixel_index2 == 4942 || pixel_index2 == 4947 || pixel_index2 == 4957 || pixel_index2 == 4964 || pixel_index2 == 4967 || pixel_index2 == 4969 || pixel_index2 == 4976 || pixel_index2 == 4978 || pixel_index2 == 4983 || pixel_index2 == 5031 || pixel_index2 == 5061 || pixel_index2 == 5221 || pixel_index2 == 5251 || ((pixel_index2 >= 5268) && (pixel_index2 <= 5270)) || pixel_index2 == 5316 || pixel_index2 == 5346 || pixel_index2 == 5367 || pixel_index2 == 5504 || pixel_index2 == 5521 || pixel_index2 == 5547 || pixel_index2 == 5550 || pixel_index2 == 5557 || ((pixel_index2 >= 5576) && (pixel_index2 <= 5579)) || ((pixel_index2 >= 5582) && (pixel_index2 <= 5583)) || ((pixel_index2 >= 5597) && (pixel_index2 <= 5599)) || ((pixel_index2 >= 5606) && (pixel_index2 <= 5607)) || ((pixel_index2 >= 5614) && (pixel_index2 <= 5616)) || ((pixel_index2 >= 5625) && (pixel_index2 <= 5628)) || ((pixel_index2 >= 5631) && (pixel_index2 <= 5632)) || ((pixel_index2 >= 5636) && (pixel_index2 <= 5637)) || ((pixel_index2 >= 5644) && (pixel_index2 <= 5645)) || (pixel_index2 >= 5650) && (pixel_index2 <= 5652)) oled_data2 = 16'b0101001010000000;
                    else if (pixel_index2 == 4909 || pixel_index2 == 4914 || ((pixel_index2 >= 4917) && (pixel_index2 <= 4922)) || ((pixel_index2 >= 4926) && (pixel_index2 <= 4929)) || ((pixel_index2 >= 4932) && (pixel_index2 <= 4933)) || pixel_index2 == 4936 || pixel_index2 == 4940 || ((pixel_index2 >= 4943) && (pixel_index2 <= 4946)) || pixel_index2 == 4958 || ((pixel_index2 >= 4962) && (pixel_index2 <= 4963)) || pixel_index2 == 4966 || ((pixel_index2 >= 4970) && (pixel_index2 <= 4975)) || ((pixel_index2 >= 4979) && (pixel_index2 <= 4982)) || ((pixel_index2 >= 5004) && (pixel_index2 <= 5005)) || ((pixel_index2 >= 5009) && (pixel_index2 <= 5010)) || ((pixel_index2 >= 5012) && (pixel_index2 <= 5019)) || ((pixel_index2 >= 5021) && (pixel_index2 <= 5026)) || ((pixel_index2 >= 5028) && (pixel_index2 <= 5030)) || ((pixel_index2 >= 5032) && (pixel_index2 <= 5033)) || ((pixel_index2 >= 5035) && (pixel_index2 <= 5036)) || ((pixel_index2 >= 5038) && (pixel_index2 <= 5043)) || ((pixel_index2 >= 5053) && (pixel_index2 <= 5054)) || ((pixel_index2 >= 5058) && (pixel_index2 <= 5060)) || ((pixel_index2 >= 5062) && (pixel_index2 <= 5063)) || ((pixel_index2 >= 5065) && (pixel_index2 <= 5072)) || ((pixel_index2 >= 5074) && (pixel_index2 <= 5079)) || ((pixel_index2 >= 5100) && (pixel_index2 <= 5101)) || ((pixel_index2 >= 5105) && (pixel_index2 <= 5106)) || ((pixel_index2 >= 5108) && (pixel_index2 <= 5110)) || ((pixel_index2 >= 5113) && (pixel_index2 <= 5115)) || ((pixel_index2 >= 5120) && (pixel_index2 <= 5122)) || ((pixel_index2 >= 5125) && (pixel_index2 <= 5129)) || ((pixel_index2 >= 5131) && (pixel_index2 <= 5132)) || ((pixel_index2 >= 5137) && (pixel_index2 <= 5139)) || ((pixel_index2 >= 5149) && (pixel_index2 <= 5150)) || ((pixel_index2 >= 5155) && (pixel_index2 <= 5159)) || ((pixel_index2 >= 5161) && (pixel_index2 <= 5163)) || ((pixel_index2 >= 5166) && (pixel_index2 <= 5168)) || ((pixel_index2 >= 5170) && (pixel_index2 <= 5172)) || ((pixel_index2 >= 5196) && (pixel_index2 <= 5197)) || ((pixel_index2 >= 5201) && (pixel_index2 <= 5202)) || ((pixel_index2 >= 5204) && (pixel_index2 <= 5205)) || ((pixel_index2 >= 5210) && (pixel_index2 <= 5211)) || ((pixel_index2 >= 5217) && (pixel_index2 <= 5218)) || ((pixel_index2 >= 5222) && (pixel_index2 <= 5225)) || ((pixel_index2 >= 5227) && (pixel_index2 <= 5228)) || ((pixel_index2 >= 5234) && (pixel_index2 <= 5235)) || ((pixel_index2 >= 5245) && (pixel_index2 <= 5246)) || ((pixel_index2 >= 5252) && (pixel_index2 <= 5255)) || ((pixel_index2 >= 5257) && (pixel_index2 <= 5258)) || ((pixel_index2 >= 5263) && (pixel_index2 <= 5264)) || ((pixel_index2 >= 5266) && (pixel_index2 <= 5267)) || ((pixel_index2 >= 5292) && (pixel_index2 <= 5293)) || ((pixel_index2 >= 5297) && (pixel_index2 <= 5298)) || ((pixel_index2 >= 5300) && (pixel_index2 <= 5301)) || ((pixel_index2 >= 5306) && (pixel_index2 <= 5307)) || ((pixel_index2 >= 5313) && (pixel_index2 <= 5314)) || ((pixel_index2 >= 5317) && (pixel_index2 <= 5321)) || ((pixel_index2 >= 5323) && (pixel_index2 <= 5324)) || ((pixel_index2 >= 5330) && (pixel_index2 <= 5331)) || ((pixel_index2 >= 5341) && (pixel_index2 <= 5342)) || ((pixel_index2 >= 5347) && (pixel_index2 <= 5351)) || ((pixel_index2 >= 5353) && (pixel_index2 <= 5354)) || ((pixel_index2 >= 5359) && (pixel_index2 <= 5360)) || ((pixel_index2 >= 5362) && (pixel_index2 <= 5366)) || ((pixel_index2 >= 5388) && (pixel_index2 <= 5389)) || ((pixel_index2 >= 5393) && (pixel_index2 <= 5394)) || ((pixel_index2 >= 5396) && (pixel_index2 <= 5397)) || ((pixel_index2 >= 5402) && (pixel_index2 <= 5403)) || ((pixel_index2 >= 5409) && (pixel_index2 <= 5410)) || ((pixel_index2 >= 5412) && (pixel_index2 <= 5414)) || ((pixel_index2 >= 5416) && (pixel_index2 <= 5417)) || ((pixel_index2 >= 5419) && (pixel_index2 <= 5420)) || ((pixel_index2 >= 5426) && (pixel_index2 <= 5427)) || ((pixel_index2 >= 5437) && (pixel_index2 <= 5438)) || ((pixel_index2 >= 5442) && (pixel_index2 <= 5444)) || ((pixel_index2 >= 5446) && (pixel_index2 <= 5447)) || ((pixel_index2 >= 5449) && (pixel_index2 <= 5450)) || ((pixel_index2 >= 5455) && (pixel_index2 <= 5456)) || ((pixel_index2 >= 5459) && (pixel_index2 <= 5463)) || ((pixel_index2 >= 5484) && (pixel_index2 <= 5485)) || ((pixel_index2 >= 5489) && (pixel_index2 <= 5490)) || ((pixel_index2 >= 5492) && (pixel_index2 <= 5493)) || ((pixel_index2 >= 5498) && (pixel_index2 <= 5499)) || ((pixel_index2 >= 5505) && (pixel_index2 <= 5506)) || ((pixel_index2 >= 5508) && (pixel_index2 <= 5509)) || ((pixel_index2 >= 5512) && (pixel_index2 <= 5513)) || ((pixel_index2 >= 5515) && (pixel_index2 <= 5516)) || ((pixel_index2 >= 5522) && (pixel_index2 <= 5523)) || ((pixel_index2 >= 5533) && (pixel_index2 <= 5534)) || ((pixel_index2 >= 5538) && (pixel_index2 <= 5539)) || ((pixel_index2 >= 5542) && (pixel_index2 <= 5543)) || ((pixel_index2 >= 5545) && (pixel_index2 <= 5546)) || ((pixel_index2 >= 5551) && (pixel_index2 <= 5552)) || ((pixel_index2 >= 5558) && (pixel_index2 <= 5559)) || ((pixel_index2 >= 5580) && (pixel_index2 <= 5581)) || ((pixel_index2 >= 5585) && (pixel_index2 <= 5586)) || ((pixel_index2 >= 5588) && (pixel_index2 <= 5589)) || ((pixel_index2 >= 5594) && (pixel_index2 <= 5595)) || ((pixel_index2 >= 5600) && (pixel_index2 <= 5602)) || ((pixel_index2 >= 5604) && (pixel_index2 <= 5605)) || ((pixel_index2 >= 5608) && (pixel_index2 <= 5609)) || ((pixel_index2 >= 5611) && (pixel_index2 <= 5612)) || ((pixel_index2 >= 5617) && (pixel_index2 <= 5619)) || ((pixel_index2 >= 5629) && (pixel_index2 <= 5630)) || ((pixel_index2 >= 5634) && (pixel_index2 <= 5635)) || ((pixel_index2 >= 5638) && (pixel_index2 <= 5639)) || ((pixel_index2 >= 5641) && (pixel_index2 <= 5643)) || ((pixel_index2 >= 5646) && (pixel_index2 <= 5648)) || ((pixel_index2 >= 5653) && (pixel_index2 <= 5655)) || ((pixel_index2 >= 5672) && (pixel_index2 <= 5679)) || ((pixel_index2 >= 5681) && (pixel_index2 <= 5682)) || ((pixel_index2 >= 5684) && (pixel_index2 <= 5685)) || ((pixel_index2 >= 5690) && (pixel_index2 <= 5691)) || ((pixel_index2 >= 5693) && (pixel_index2 <= 5698)) || ((pixel_index2 >= 5700) && (pixel_index2 <= 5705)) || ((pixel_index2 >= 5707) && (pixel_index2 <= 5708)) || ((pixel_index2 >= 5710) && (pixel_index2 <= 5715)) || ((pixel_index2 >= 5721) && (pixel_index2 <= 5728)) || ((pixel_index2 >= 5730) && (pixel_index2 <= 5735)) || ((pixel_index2 >= 5737) && (pixel_index2 <= 5744)) || ((pixel_index2 >= 5746) && (pixel_index2 <= 5751)) || ((pixel_index2 >= 5769) && (pixel_index2 <= 5774)) || pixel_index2 == 5777 || pixel_index2 == 5781 || pixel_index2 == 5786 || ((pixel_index2 >= 5790) && (pixel_index2 <= 5793)) || ((pixel_index2 >= 5797) && (pixel_index2 <= 5800)) || pixel_index2 == 5803 || ((pixel_index2 >= 5807) && (pixel_index2 <= 5810)) || ((pixel_index2 >= 5818) && (pixel_index2 <= 5823)) || ((pixel_index2 >= 5827) && (pixel_index2 <= 5830)) || ((pixel_index2 >= 5834) && (pixel_index2 <= 5839)) || (pixel_index2 >= 5843) && (pixel_index2 <= 5846)) oled_data2 = 16'b1111010100010100;
                    else oled_data2 = 0;
                end
                2: begin
                    if (pixel_index2 == 97 || pixel_index2 == 99 || pixel_index2 == 101 || ((pixel_index2 >= 103) && (pixel_index2 <= 104)) || ((pixel_index2 >= 106) && (pixel_index2 <= 109)) || pixel_index2 == 111 || ((pixel_index2 >= 113) && (pixel_index2 <= 114)) || ((pixel_index2 >= 118) && (pixel_index2 <= 120)) || pixel_index2 == 195 || pixel_index2 == 197 || ((pixel_index2 >= 199) && (pixel_index2 <= 200)) || pixel_index2 == 202 || ((pixel_index2 >= 204) && (pixel_index2 <= 205)) || pixel_index2 == 207 || ((pixel_index2 >= 209) && (pixel_index2 <= 210)) || pixel_index2 == 213 || pixel_index2 == 289 || ((pixel_index2 >= 291) && (pixel_index2 <= 296)) || pixel_index2 == 298 || ((pixel_index2 >= 300) && (pixel_index2 <= 301)) || pixel_index2 == 303 || ((pixel_index2 >= 305) && (pixel_index2 <= 306)) || ((pixel_index2 >= 310) && (pixel_index2 <= 312)) || pixel_index2 == 385 || ((pixel_index2 >= 387) && (pixel_index2 <= 392)) || pixel_index2 == 394 || ((pixel_index2 >= 396) && (pixel_index2 <= 397)) || ((pixel_index2 >= 399) && (pixel_index2 <= 402)) || pixel_index2 == 408 || ((pixel_index2 >= 501) && (pixel_index2 <= 504)) || ((pixel_index2 >= 674) && (pixel_index2 <= 675)) || ((pixel_index2 >= 678) && (pixel_index2 <= 681)) || ((pixel_index2 >= 685) && (pixel_index2 <= 686)) || pixel_index2 == 688 || ((pixel_index2 >= 690) && (pixel_index2 <= 691)) || ((pixel_index2 >= 693) && (pixel_index2 <= 696)) || ((pixel_index2 >= 770) && (pixel_index2 <= 771)) || pixel_index2 == 774 || ((pixel_index2 >= 776) && (pixel_index2 <= 777)) || ((pixel_index2 >= 779) && (pixel_index2 <= 782)) || pixel_index2 == 784 || ((pixel_index2 >= 786) && (pixel_index2 <= 787)) || ((pixel_index2 >= 790) && (pixel_index2 <= 791)) || ((pixel_index2 >= 866) && (pixel_index2 <= 867)) || pixel_index2 == 870 || ((pixel_index2 >= 872) && (pixel_index2 <= 873)) || pixel_index2 == 875 || ((pixel_index2 >= 877) && (pixel_index2 <= 878)) || pixel_index2 == 880 || ((pixel_index2 >= 882) && (pixel_index2 <= 883)) || ((pixel_index2 >= 886) && (pixel_index2 <= 887)) || ((pixel_index2 >= 895) && (pixel_index2 <= 896)) || ((pixel_index2 >= 899) && (pixel_index2 <= 900)) || ((pixel_index2 >= 903) && (pixel_index2 <= 904)) || ((pixel_index2 >= 907) && (pixel_index2 <= 908)) || ((pixel_index2 >= 911) && (pixel_index2 <= 912)) || ((pixel_index2 >= 915) && (pixel_index2 <= 916)) || ((pixel_index2 >= 919) && (pixel_index2 <= 920)) || ((pixel_index2 >= 923) && (pixel_index2 <= 924)) || ((pixel_index2 >= 927) && (pixel_index2 <= 928)) || ((pixel_index2 >= 931) && (pixel_index2 <= 932)) || ((pixel_index2 >= 935) && (pixel_index2 <= 936)) || ((pixel_index2 >= 939) && (pixel_index2 <= 940)) || ((pixel_index2 >= 943) && (pixel_index2 <= 944)) || ((pixel_index2 >= 947) && (pixel_index2 <= 948)) || ((pixel_index2 >= 951) && (pixel_index2 <= 952)) || ((pixel_index2 >= 955) && (pixel_index2 <= 956)) || ((pixel_index2 >= 961) && (pixel_index2 <= 964)) || pixel_index2 == 966 || ((pixel_index2 >= 968) && (pixel_index2 <= 969)) || ((pixel_index2 >= 971) && (pixel_index2 <= 974)) || ((pixel_index2 >= 976) && (pixel_index2 <= 979)) || ((pixel_index2 >= 981) && (pixel_index2 <= 984)) || pixel_index2 == 1155 || ((pixel_index2 >= 1159) && (pixel_index2 <= 1161)) || pixel_index2 == 1163 || ((pixel_index2 >= 1165) && (pixel_index2 <= 1166)) || pixel_index2 == 1168 || ((pixel_index2 >= 1170) && (pixel_index2 <= 1171)) || pixel_index2 == 1173 || ((pixel_index2 >= 1175) && (pixel_index2 <= 1176)) || pixel_index2 == 1254 || ((pixel_index2 >= 1256) && (pixel_index2 <= 1257)) || pixel_index2 == 1259 || ((pixel_index2 >= 1261) && (pixel_index2 <= 1262)) || ((pixel_index2 >= 1264) && (pixel_index2 <= 1267)) || ((pixel_index2 >= 1270) && (pixel_index2 <= 1272)) || pixel_index2 == 1350 || ((pixel_index2 >= 1352) && (pixel_index2 <= 1353)) || pixel_index2 == 1355 || ((pixel_index2 >= 1357) && (pixel_index2 <= 1358)) || pixel_index2 == 1360 || ((pixel_index2 >= 1362) && (pixel_index2 <= 1363)) || pixel_index2 == 1365 || ((pixel_index2 >= 1367) && (pixel_index2 <= 1368)) || ((pixel_index2 >= 1447) && (pixel_index2 <= 1449)) || ((pixel_index2 >= 1451) && (pixel_index2 <= 1454)) || ((pixel_index2 >= 1456) && (pixel_index2 <= 1459)) || ((pixel_index2 >= 1461) && (pixel_index2 <= 1464)) || ((pixel_index2 >= 1637) && (pixel_index2 <= 1638)) || ((pixel_index2 >= 1641) && (pixel_index2 <= 1644)) || ((pixel_index2 >= 1646) && (pixel_index2 <= 1649)) || ((pixel_index2 >= 1652) && (pixel_index2 <= 1654)) || pixel_index2 == 1732 || pixel_index2 == 1735 || pixel_index2 == 1740 || pixel_index2 == 1745 || pixel_index2 == 1747 || pixel_index2 == 1831 || pixel_index2 == 1836 || ((pixel_index2 >= 1839) && (pixel_index2 <= 1841)) || ((pixel_index2 >= 1844) && (pixel_index2 <= 1845)) || pixel_index2 == 1924 || pixel_index2 == 1927 || pixel_index2 == 1932 || pixel_index2 == 1937 || pixel_index2 == 1942 || ((pixel_index2 >= 2021) && (pixel_index2 <= 2022)) || pixel_index2 == 2028 || ((pixel_index2 >= 2030) && (pixel_index2 <= 2033)) || ((pixel_index2 >= 2035) && (pixel_index2 <= 2037)) || pixel_index2 == 2213 || pixel_index2 == 2216 || ((pixel_index2 >= 2219) && (pixel_index2 <= 2221)) || pixel_index2 == 2223 || pixel_index2 == 2226 || ((pixel_index2 >= 2228) && (pixel_index2 <= 2230)) || pixel_index2 == 2310 || pixel_index2 == 2312 || pixel_index2 == 2314 || pixel_index2 == 2319 || pixel_index2 == 2322 || pixel_index2 == 2325 || ((pixel_index2 >= 2406) && (pixel_index2 <= 2408)) || ((pixel_index2 >= 2411) && (pixel_index2 <= 2412)) || ((pixel_index2 >= 2415) && (pixel_index2 <= 2416)) || pixel_index2 == 2418 || pixel_index2 == 2421 || pixel_index2 == 2501 || pixel_index2 == 2504 || pixel_index2 == 2509 || pixel_index2 == 2511 || ((pixel_index2 >= 2513) && (pixel_index2 <= 2514)) || pixel_index2 == 2517 || ((pixel_index2 >= 2598) && (pixel_index2 <= 2600)) || ((pixel_index2 >= 2602) && (pixel_index2 <= 2604)) || pixel_index2 == 2607 || pixel_index2 == 2610 || ((pixel_index2 >= 2612) && (pixel_index2 <= 2614)) || pixel_index2 == 2788 || pixel_index2 == 2791 || ((pixel_index2 >= 2794) && (pixel_index2 <= 2795)) || ((pixel_index2 >= 2799) && (pixel_index2 <= 2800)) || ((pixel_index2 >= 2804) && (pixel_index2 <= 2805)) || pixel_index2 == 2885 || pixel_index2 == 2887 || pixel_index2 == 2889 || pixel_index2 == 2892 || pixel_index2 == 2894 || pixel_index2 == 2897 || pixel_index2 == 2899 || pixel_index2 == 2902 || ((pixel_index2 >= 2982) && (pixel_index2 <= 2983)) || pixel_index2 == 2988 || pixel_index2 == 2990 || pixel_index2 == 2993 || pixel_index2 == 2998 || pixel_index2 == 3077 || pixel_index2 == 3079 || pixel_index2 == 3081 || pixel_index2 == 3084 || pixel_index2 == 3086 || pixel_index2 == 3089 || pixel_index2 == 3091 || pixel_index2 == 3094 || ((pixel_index2 >= 3133) && (pixel_index2 <= 3134)) || pixel_index2 == 3172 || pixel_index2 == 3175 || ((pixel_index2 >= 3178) && (pixel_index2 <= 3179)) || ((pixel_index2 >= 3183) && (pixel_index2 <= 3184)) || ((pixel_index2 >= 3188) && (pixel_index2 <= 3189)) || pixel_index2 == 3228 || pixel_index2 == 3327 || ((pixel_index2 >= 3364) && (pixel_index2 <= 3367)) || ((pixel_index2 >= 3370) && (pixel_index2 <= 3372)) || ((pixel_index2 >= 3375) && (pixel_index2 <= 3376)) || ((pixel_index2 >= 3380) && (pixel_index2 <= 3382)) || pixel_index2 == 3463 || pixel_index2 == 3465 || pixel_index2 == 3468 || pixel_index2 == 3470 || pixel_index2 == 3473 || pixel_index2 == 3475 || pixel_index2 == 3478 || pixel_index2 == 3559 || ((pixel_index2 >= 3562) && (pixel_index2 <= 3564)) || pixel_index2 == 3566 || pixel_index2 == 3569 || ((pixel_index2 >= 3572) && (pixel_index2 <= 3574)) || ((pixel_index2 >= 3630) && (pixel_index2 <= 3631)) || pixel_index2 == 3655 || pixel_index2 == 3657 || pixel_index2 == 3660 || pixel_index2 == 3662 || pixel_index2 == 3665 || pixel_index2 == 3667 || pixel_index2 == 3670 || pixel_index2 == 3751 || ((pixel_index2 >= 3754) && (pixel_index2 <= 3756)) || pixel_index2 == 3758 || pixel_index2 == 3761 || ((pixel_index2 >= 3764) && (pixel_index2 <= 3766)) || ((pixel_index2 >= 4008) && (pixel_index2 <= 4009)) || ((pixel_index2 >= 4012) && (pixel_index2 <= 4015)) || ((pixel_index2 >= 4017) && (pixel_index2 <= 4020)) || ((pixel_index2 >= 4022) && (pixel_index2 <= 4025)) || pixel_index2 == 4027 || ((pixel_index2 >= 4029) && (pixel_index2 <= 4030)) || ((pixel_index2 >= 4104) && (pixel_index2 <= 4105)) || ((pixel_index2 >= 4110) && (pixel_index2 <= 4111)) || ((pixel_index2 >= 4113) && (pixel_index2 <= 4114)) || ((pixel_index2 >= 4120) && (pixel_index2 <= 4121)) || ((pixel_index2 >= 4124) && (pixel_index2 <= 4126)) || ((pixel_index2 >= 4200) && (pixel_index2 <= 4201)) || ((pixel_index2 >= 4204) && (pixel_index2 <= 4205)) || pixel_index2 == 4207 || ((pixel_index2 >= 4210) && (pixel_index2 <= 4212)) || ((pixel_index2 >= 4214) && (pixel_index2 <= 4215)) || pixel_index2 == 4217 || pixel_index2 == 4219 || ((pixel_index2 >= 4221) && (pixel_index2 <= 4222)) || ((pixel_index2 >= 4295) && (pixel_index2 <= 4298)) || ((pixel_index2 >= 4300) && (pixel_index2 <= 4303)) || ((pixel_index2 >= 4305) && (pixel_index2 <= 4307)) || ((pixel_index2 >= 4310) && (pixel_index2 <= 4313)) || ((pixel_index2 >= 4315) && (pixel_index2 <= 4318)) || pixel_index2 == 4802 || pixel_index2 == 4893 || pixel_index2 == 5762 || pixel_index2 == 5853) oled_data2 = 16'b1111011110011110;
                    else if (((pixel_index2 >= 124) && (pixel_index2 <= 190)) || ((pixel_index2 >= 220) && (pixel_index2 <= 221)) || pixel_index2 == 225 || pixel_index2 == 229 || pixel_index2 == 233 || pixel_index2 == 237 || pixel_index2 == 241 || pixel_index2 == 245 || pixel_index2 == 249 || pixel_index2 == 253 || pixel_index2 == 257 || pixel_index2 == 261 || pixel_index2 == 265 || pixel_index2 == 269 || pixel_index2 == 273 || pixel_index2 == 277 || pixel_index2 == 281 || ((pixel_index2 >= 285) && (pixel_index2 <= 286)) || ((pixel_index2 >= 316) && (pixel_index2 <= 317)) || pixel_index2 == 321 || pixel_index2 == 325 || pixel_index2 == 329 || pixel_index2 == 333 || pixel_index2 == 337 || pixel_index2 == 341 || pixel_index2 == 345 || pixel_index2 == 349 || pixel_index2 == 353 || pixel_index2 == 357 || pixel_index2 == 361 || pixel_index2 == 365 || pixel_index2 == 369 || pixel_index2 == 373 || pixel_index2 == 377 || ((pixel_index2 >= 381) && (pixel_index2 <= 382)) || ((pixel_index2 >= 412) && (pixel_index2 <= 413)) || pixel_index2 == 417 || pixel_index2 == 421 || pixel_index2 == 425 || pixel_index2 == 429 || pixel_index2 == 433 || pixel_index2 == 437 || pixel_index2 == 441 || pixel_index2 == 445 || pixel_index2 == 449 || pixel_index2 == 453 || pixel_index2 == 457 || pixel_index2 == 461 || pixel_index2 == 465 || pixel_index2 == 469 || pixel_index2 == 473 || ((pixel_index2 >= 477) && (pixel_index2 <= 478)) || ((pixel_index2 >= 508) && (pixel_index2 <= 509)) || pixel_index2 == 513 || pixel_index2 == 517 || pixel_index2 == 521 || pixel_index2 == 525 || pixel_index2 == 529 || pixel_index2 == 533 || pixel_index2 == 537 || pixel_index2 == 541 || pixel_index2 == 545 || pixel_index2 == 549 || pixel_index2 == 553 || pixel_index2 == 557 || pixel_index2 == 561 || pixel_index2 == 565 || pixel_index2 == 569 || ((pixel_index2 >= 573) && (pixel_index2 <= 574)) || ((pixel_index2 >= 604) && (pixel_index2 <= 605)) || pixel_index2 == 609 || pixel_index2 == 613 || pixel_index2 == 617 || pixel_index2 == 621 || pixel_index2 == 625 || pixel_index2 == 629 || pixel_index2 == 633 || pixel_index2 == 637 || pixel_index2 == 641 || pixel_index2 == 645 || pixel_index2 == 649 || pixel_index2 == 653 || pixel_index2 == 657 || pixel_index2 == 661 || pixel_index2 == 665 || ((pixel_index2 >= 669) && (pixel_index2 <= 670)) || ((pixel_index2 >= 700) && (pixel_index2 <= 701)) || pixel_index2 == 705 || pixel_index2 == 709 || pixel_index2 == 713 || pixel_index2 == 717 || pixel_index2 == 721 || pixel_index2 == 725 || pixel_index2 == 729 || pixel_index2 == 733 || pixel_index2 == 737 || pixel_index2 == 741 || pixel_index2 == 745 || pixel_index2 == 749 || pixel_index2 == 753 || pixel_index2 == 757 || pixel_index2 == 761 || ((pixel_index2 >= 765) && (pixel_index2 <= 766)) || ((pixel_index2 >= 796) && (pixel_index2 <= 862)) || ((pixel_index2 >= 892) && (pixel_index2 <= 894)) || ((pixel_index2 >= 897) && (pixel_index2 <= 898)) || ((pixel_index2 >= 901) && (pixel_index2 <= 902)) || ((pixel_index2 >= 905) && (pixel_index2 <= 906)) || ((pixel_index2 >= 909) && (pixel_index2 <= 910)) || ((pixel_index2 >= 913) && (pixel_index2 <= 914)) || ((pixel_index2 >= 917) && (pixel_index2 <= 918)) || ((pixel_index2 >= 921) && (pixel_index2 <= 922)) || ((pixel_index2 >= 925) && (pixel_index2 <= 926)) || ((pixel_index2 >= 929) && (pixel_index2 <= 930)) || ((pixel_index2 >= 933) && (pixel_index2 <= 934)) || ((pixel_index2 >= 937) && (pixel_index2 <= 938)) || ((pixel_index2 >= 941) && (pixel_index2 <= 942)) || ((pixel_index2 >= 945) && (pixel_index2 <= 946)) || ((pixel_index2 >= 949) && (pixel_index2 <= 950)) || ((pixel_index2 >= 953) && (pixel_index2 <= 954)) || ((pixel_index2 >= 957) && (pixel_index2 <= 958)) || ((pixel_index2 >= 988) && (pixel_index2 <= 1054)) || ((pixel_index2 >= 1084) && (pixel_index2 <= 1085)) || ((pixel_index2 >= 1087) && (pixel_index2 <= 1089)) || ((pixel_index2 >= 1091) && (pixel_index2 <= 1093)) || ((pixel_index2 >= 1095) && (pixel_index2 <= 1097)) || ((pixel_index2 >= 1099) && (pixel_index2 <= 1101)) || ((pixel_index2 >= 1103) && (pixel_index2 <= 1105)) || ((pixel_index2 >= 1107) && (pixel_index2 <= 1109)) || ((pixel_index2 >= 1111) && (pixel_index2 <= 1113)) || ((pixel_index2 >= 1115) && (pixel_index2 <= 1117)) || ((pixel_index2 >= 1119) && (pixel_index2 <= 1121)) || ((pixel_index2 >= 1123) && (pixel_index2 <= 1125)) || ((pixel_index2 >= 1127) && (pixel_index2 <= 1129)) || ((pixel_index2 >= 1131) && (pixel_index2 <= 1133)) || ((pixel_index2 >= 1135) && (pixel_index2 <= 1137)) || ((pixel_index2 >= 1139) && (pixel_index2 <= 1141)) || ((pixel_index2 >= 1143) && (pixel_index2 <= 1145)) || ((pixel_index2 >= 1147) && (pixel_index2 <= 1150)) || ((pixel_index2 >= 1182) && (pixel_index2 <= 1219)) || ((pixel_index2 >= 1240) && (pixel_index2 <= 1244)) || ((pixel_index2 >= 1278) && (pixel_index2 <= 1280)) || ((pixel_index2 >= 1283) && (pixel_index2 <= 1286)) || ((pixel_index2 >= 1290) && (pixel_index2 <= 1291)) || ((pixel_index2 >= 1293) && (pixel_index2 <= 1294)) || ((pixel_index2 >= 1314) && (pixel_index2 <= 1315)) || ((pixel_index2 >= 1336) && (pixel_index2 <= 1340)) || ((pixel_index2 >= 1374) && (pixel_index2 <= 1376)) || ((pixel_index2 >= 1378) && (pixel_index2 <= 1382)) || ((pixel_index2 >= 1386) && (pixel_index2 <= 1390)) || ((pixel_index2 >= 1410) && (pixel_index2 <= 1411)) || ((pixel_index2 >= 1432) && (pixel_index2 <= 1436)) || ((pixel_index2 >= 1470) && (pixel_index2 <= 1478)) || ((pixel_index2 >= 1482) && (pixel_index2 <= 1486)) || ((pixel_index2 >= 1506) && (pixel_index2 <= 1507)) || ((pixel_index2 >= 1528) && (pixel_index2 <= 1532)) || ((pixel_index2 >= 1566) && (pixel_index2 <= 1573)) || ((pixel_index2 >= 1579) && (pixel_index2 <= 1603)) || ((pixel_index2 >= 1624) && (pixel_index2 <= 1628)) || ((pixel_index2 >= 1662) && (pixel_index2 <= 1666)) || ((pixel_index2 >= 1678) && (pixel_index2 <= 1696)) || ((pixel_index2 >= 1698) && (pixel_index2 <= 1699)) || ((pixel_index2 >= 1720) && (pixel_index2 <= 1724)) || ((pixel_index2 >= 1758) && (pixel_index2 <= 1762)) || ((pixel_index2 >= 1774) && (pixel_index2 <= 1775)) || ((pixel_index2 >= 1777) && (pixel_index2 <= 1789)) || pixel_index2 == 1792 || ((pixel_index2 >= 1794) && (pixel_index2 <= 1795)) || pixel_index2 == 1816 || ((pixel_index2 >= 1818) && (pixel_index2 <= 1820)) || ((pixel_index2 >= 1854) && (pixel_index2 <= 1858)) || pixel_index2 == 1870 || ((pixel_index2 >= 1872) && (pixel_index2 <= 1878)) || ((pixel_index2 >= 1882) && (pixel_index2 <= 1888)) || ((pixel_index2 >= 1892) && (pixel_index2 <= 1913)) || ((pixel_index2 >= 1915) && (pixel_index2 <= 1916)) || ((pixel_index2 >= 1948) && (pixel_index2 <= 1957)) || ((pixel_index2 >= 1963) && (pixel_index2 <= 1973)) || pixel_index2 == 1988 || pixel_index2 == 1991 || ((pixel_index2 >= 1993) && (pixel_index2 <= 1994)) || pixel_index2 == 1996 || ((pixel_index2 >= 2000) && (pixel_index2 <= 2001)) || pixel_index2 == 2008 || ((pixel_index2 >= 2011) && (pixel_index2 <= 2014)) || ((pixel_index2 >= 2044) && (pixel_index2 <= 2046)) || ((pixel_index2 >= 2048) && (pixel_index2 <= 2054)) || ((pixel_index2 >= 2058) && (pixel_index2 <= 2069)) || ((pixel_index2 >= 2084) && (pixel_index2 <= 2085)) || pixel_index2 == 2089 || ((pixel_index2 >= 2091) && (pixel_index2 <= 2093)) || ((pixel_index2 >= 2095) && (pixel_index2 <= 2096)) || ((pixel_index2 >= 2104) && (pixel_index2 <= 2105)) || ((pixel_index2 >= 2107) && (pixel_index2 <= 2110)) || pixel_index2 == 2140 || pixel_index2 == 2142 || ((pixel_index2 >= 2144) && (pixel_index2 <= 2150)) || pixel_index2 == 2154 || ((pixel_index2 >= 2157) && (pixel_index2 <= 2168)) || pixel_index2 == 2178 || ((pixel_index2 >= 2180) && (pixel_index2 <= 2184)) || pixel_index2 == 2188 || ((pixel_index2 >= 2190) && (pixel_index2 <= 2192)) || ((pixel_index2 >= 2195) && (pixel_index2 <= 2197)) || ((pixel_index2 >= 2200) && (pixel_index2 <= 2206)) || ((pixel_index2 >= 2236) && (pixel_index2 <= 2238)) || ((pixel_index2 >= 2245) && (pixel_index2 <= 2246)) || pixel_index2 == 2250 || ((pixel_index2 >= 2252) && (pixel_index2 <= 2264)) || ((pixel_index2 >= 2274) && (pixel_index2 <= 2288)) || ((pixel_index2 >= 2291) && (pixel_index2 <= 2293)) || ((pixel_index2 >= 2296) && (pixel_index2 <= 2302)) || ((pixel_index2 >= 2332) && (pixel_index2 <= 2334)) || ((pixel_index2 >= 2341) && (pixel_index2 <= 2355)) || ((pixel_index2 >= 2374) && (pixel_index2 <= 2384)) || ((pixel_index2 >= 2392) && (pixel_index2 <= 2398)) || ((pixel_index2 >= 2428) && (pixel_index2 <= 2437)) || ((pixel_index2 >= 2443) && (pixel_index2 <= 2451)) || ((pixel_index2 >= 2470) && (pixel_index2 <= 2480)) || ((pixel_index2 >= 2487) && (pixel_index2 <= 2494)) || ((pixel_index2 >= 2526) && (pixel_index2 <= 2532)) || ((pixel_index2 >= 2540) && (pixel_index2 <= 2547)) || pixel_index2 == 2566 || ((pixel_index2 >= 2580) && (pixel_index2 <= 2588)) || ((pixel_index2 >= 2622) && (pixel_index2 <= 2626)) || pixel_index2 == 2636 || ((pixel_index2 >= 2639) && (pixel_index2 <= 2644)) || ((pixel_index2 >= 2647) && (pixel_index2 <= 2648)) || pixel_index2 == 2659 || ((pixel_index2 >= 2661) && (pixel_index2 <= 2662)) || ((pixel_index2 >= 2676) && (pixel_index2 <= 2684)) || ((pixel_index2 >= 2718) && (pixel_index2 <= 2721)) || pixel_index2 == 2732 || ((pixel_index2 >= 2735) && (pixel_index2 <= 2742)) || ((pixel_index2 >= 2756) && (pixel_index2 <= 2758)) || ((pixel_index2 >= 2772) && (pixel_index2 <= 2780)) || ((pixel_index2 >= 2814) && (pixel_index2 <= 2817)) || pixel_index2 == 2828 || ((pixel_index2 >= 2831) && (pixel_index2 <= 2838)) || ((pixel_index2 >= 2842) && (pixel_index2 <= 2848)) || ((pixel_index2 >= 2852) && (pixel_index2 <= 2859)) || ((pixel_index2 >= 2866) && (pixel_index2 <= 2876)) || ((pixel_index2 >= 2910) && (pixel_index2 <= 2913)) || pixel_index2 == 2924 || ((pixel_index2 >= 2927) && (pixel_index2 <= 2935)) || ((pixel_index2 >= 2938) && (pixel_index2 <= 2944)) || ((pixel_index2 >= 2947) && (pixel_index2 <= 2955)) || pixel_index2 == 2962 || ((pixel_index2 >= 2964) && (pixel_index2 <= 2972)) || ((pixel_index2 >= 3006) && (pixel_index2 <= 3013)) || ((pixel_index2 >= 3019) && (pixel_index2 <= 3021)) || ((pixel_index2 >= 3023) && (pixel_index2 <= 3032)) || ((pixel_index2 >= 3042) && (pixel_index2 <= 3051)) || ((pixel_index2 >= 3058) && (pixel_index2 <= 3060)) || pixel_index2 == 3063 || ((pixel_index2 >= 3065) && (pixel_index2 <= 3068)) || ((pixel_index2 >= 3102) && (pixel_index2 <= 3104)) || pixel_index2 == 3107 || ((pixel_index2 >= 3117) && (pixel_index2 <= 3123)) || ((pixel_index2 >= 3143) && (pixel_index2 <= 3147)) || ((pixel_index2 >= 3154) && (pixel_index2 <= 3155)) || pixel_index2 == 3159 || ((pixel_index2 >= 3161) && (pixel_index2 <= 3164)) || ((pixel_index2 >= 3198) && (pixel_index2 <= 3200)) || ((pixel_index2 >= 3202) && (pixel_index2 <= 3203)) || ((pixel_index2 >= 3213) && (pixel_index2 <= 3216)) || ((pixel_index2 >= 3218) && (pixel_index2 <= 3219)) || ((pixel_index2 >= 3239) && (pixel_index2 <= 3243)) || ((pixel_index2 >= 3250) && (pixel_index2 <= 3251)) || ((pixel_index2 >= 3255) && (pixel_index2 <= 3260)) || ((pixel_index2 >= 3292) && (pixel_index2 <= 3299)) || ((pixel_index2 >= 3309) && (pixel_index2 <= 3312)) || ((pixel_index2 >= 3314) && (pixel_index2 <= 3315)) || ((pixel_index2 >= 3335) && (pixel_index2 <= 3337)) || pixel_index2 == 3339 || ((pixel_index2 >= 3346) && (pixel_index2 <= 3347)) || ((pixel_index2 >= 3351) && (pixel_index2 <= 3352)) || ((pixel_index2 >= 3354) && (pixel_index2 <= 3358)) || ((pixel_index2 >= 3388) && (pixel_index2 <= 3393)) || pixel_index2 == 3395 || ((pixel_index2 >= 3405) && (pixel_index2 <= 3407)) || ((pixel_index2 >= 3409) && (pixel_index2 <= 3411)) || ((pixel_index2 >= 3431) && (pixel_index2 <= 3432)) || ((pixel_index2 >= 3434) && (pixel_index2 <= 3435)) || ((pixel_index2 >= 3438) && (pixel_index2 <= 3443)) || ((pixel_index2 >= 3447) && (pixel_index2 <= 3448)) || ((pixel_index2 >= 3450) && (pixel_index2 <= 3454)) || ((pixel_index2 >= 3484) && (pixel_index2 <= 3487)) || pixel_index2 == 3489 || pixel_index2 == 3491 || ((pixel_index2 >= 3501) && (pixel_index2 <= 3502)) || ((pixel_index2 >= 3505) && (pixel_index2 <= 3507)) || ((pixel_index2 >= 3527) && (pixel_index2 <= 3531)) || ((pixel_index2 >= 3538) && (pixel_index2 <= 3539)) || ((pixel_index2 >= 3543) && (pixel_index2 <= 3544)) || ((pixel_index2 >= 3546) && (pixel_index2 <= 3550)) || ((pixel_index2 >= 3580) && (pixel_index2 <= 3587)) || ((pixel_index2 >= 3597) && (pixel_index2 <= 3603)) || ((pixel_index2 >= 3623) && (pixel_index2 <= 3628)) || ((pixel_index2 >= 3633) && (pixel_index2 <= 3635)) || ((pixel_index2 >= 3639) && (pixel_index2 <= 3646)) || ((pixel_index2 >= 4620) && (pixel_index2 <= 4692)) || ((pixel_index2 >= 4707) && (pixel_index2 <= 4796)) || ((pixel_index2 >= 4803) && (pixel_index2 <= 4812)) || ((pixel_index2 >= 4814) && (pixel_index2 <= 4817)) || ((pixel_index2 >= 4819) && (pixel_index2 <= 4820)) || ((pixel_index2 >= 4827) && (pixel_index2 <= 4829)) || ((pixel_index2 >= 4834) && (pixel_index2 <= 4835)) || ((pixel_index2 >= 4838) && (pixel_index2 <= 4839)) || ((pixel_index2 >= 4841) && (pixel_index2 <= 4843)) || ((pixel_index2 >= 4845) && (pixel_index2 <= 4846)) || ((pixel_index2 >= 4851) && (pixel_index2 <= 4861)) || ((pixel_index2 >= 4863) && (pixel_index2 <= 4865)) || ((pixel_index2 >= 4868) && (pixel_index2 <= 4869)) || ((pixel_index2 >= 4871) && (pixel_index2 <= 4873)) || ((pixel_index2 >= 4880) && (pixel_index2 <= 4882)) || ((pixel_index2 >= 4887) && (pixel_index2 <= 4892)) || ((pixel_index2 >= 4899) && (pixel_index2 <= 4907)) || ((pixel_index2 >= 4910) && (pixel_index2 <= 4912)) || pixel_index2 == 4915 || pixel_index2 == 4924 || pixel_index2 == 4931 || pixel_index2 == 4935 || pixel_index2 == 4938 || pixel_index2 == 4941 || ((pixel_index2 >= 4948) && (pixel_index2 <= 4956)) || ((pixel_index2 >= 4959) && (pixel_index2 <= 4961)) || pixel_index2 == 4965 || pixel_index2 == 4968 || pixel_index2 == 4977 || ((pixel_index2 >= 4984) && (pixel_index2 <= 4988)) || ((pixel_index2 >= 4994) && (pixel_index2 <= 5003)) || ((pixel_index2 >= 5006) && (pixel_index2 <= 5008)) || pixel_index2 == 5011 || pixel_index2 == 5020 || pixel_index2 == 5027 || pixel_index2 == 5034 || pixel_index2 == 5037 || ((pixel_index2 >= 5044) && (pixel_index2 <= 5052)) || ((pixel_index2 >= 5055) && (pixel_index2 <= 5057)) || pixel_index2 == 5064 || pixel_index2 == 5073 || ((pixel_index2 >= 5080) && (pixel_index2 <= 5085)) || ((pixel_index2 >= 5090) && (pixel_index2 <= 5099)) || ((pixel_index2 >= 5102) && (pixel_index2 <= 5104)) || pixel_index2 == 5107 || ((pixel_index2 >= 5111) && (pixel_index2 <= 5112)) || ((pixel_index2 >= 5116) && (pixel_index2 <= 5119)) || ((pixel_index2 >= 5123) && (pixel_index2 <= 5124)) || pixel_index2 == 5130 || ((pixel_index2 >= 5133) && (pixel_index2 <= 5136)) || ((pixel_index2 >= 5140) && (pixel_index2 <= 5148)) || ((pixel_index2 >= 5151) && (pixel_index2 <= 5154)) || pixel_index2 == 5160 || ((pixel_index2 >= 5164) && (pixel_index2 <= 5165)) || pixel_index2 == 5169 || ((pixel_index2 >= 5173) && (pixel_index2 <= 5181)) || ((pixel_index2 >= 5186) && (pixel_index2 <= 5195)) || ((pixel_index2 >= 5198) && (pixel_index2 <= 5200)) || pixel_index2 == 5203 || ((pixel_index2 >= 5206) && (pixel_index2 <= 5209)) || ((pixel_index2 >= 5212) && (pixel_index2 <= 5216)) || ((pixel_index2 >= 5219) && (pixel_index2 <= 5220)) || pixel_index2 == 5226 || ((pixel_index2 >= 5229) && (pixel_index2 <= 5233)) || ((pixel_index2 >= 5236) && (pixel_index2 <= 5244)) || ((pixel_index2 >= 5247) && (pixel_index2 <= 5250)) || pixel_index2 == 5256 || ((pixel_index2 >= 5259) && (pixel_index2 <= 5262)) || pixel_index2 == 5265 || ((pixel_index2 >= 5271) && (pixel_index2 <= 5277)) || ((pixel_index2 >= 5282) && (pixel_index2 <= 5291)) || ((pixel_index2 >= 5294) && (pixel_index2 <= 5296)) || pixel_index2 == 5299 || ((pixel_index2 >= 5302) && (pixel_index2 <= 5305)) || ((pixel_index2 >= 5308) && (pixel_index2 <= 5312)) || pixel_index2 == 5315 || pixel_index2 == 5322 || ((pixel_index2 >= 5325) && (pixel_index2 <= 5329)) || ((pixel_index2 >= 5332) && (pixel_index2 <= 5340)) || ((pixel_index2 >= 5343) && (pixel_index2 <= 5345)) || pixel_index2 == 5352 || ((pixel_index2 >= 5355) && (pixel_index2 <= 5358)) || pixel_index2 == 5361 || ((pixel_index2 >= 5368) && (pixel_index2 <= 5373)) || ((pixel_index2 >= 5378) && (pixel_index2 <= 5387)) || ((pixel_index2 >= 5390) && (pixel_index2 <= 5392)) || pixel_index2 == 5395 || ((pixel_index2 >= 5398) && (pixel_index2 <= 5401)) || ((pixel_index2 >= 5404) && (pixel_index2 <= 5408)) || pixel_index2 == 5411 || pixel_index2 == 5415 || pixel_index2 == 5418 || ((pixel_index2 >= 5421) && (pixel_index2 <= 5425)) || ((pixel_index2 >= 5428) && (pixel_index2 <= 5436)) || ((pixel_index2 >= 5439) && (pixel_index2 <= 5441)) || pixel_index2 == 5445 || pixel_index2 == 5448 || ((pixel_index2 >= 5451) && (pixel_index2 <= 5454)) || ((pixel_index2 >= 5457) && (pixel_index2 <= 5458)) || ((pixel_index2 >= 5464) && (pixel_index2 <= 5469)) || ((pixel_index2 >= 5474) && (pixel_index2 <= 5483)) || ((pixel_index2 >= 5486) && (pixel_index2 <= 5488)) || pixel_index2 == 5491 || ((pixel_index2 >= 5494) && (pixel_index2 <= 5497)) || ((pixel_index2 >= 5500) && (pixel_index2 <= 5503)) || pixel_index2 == 5507 || ((pixel_index2 >= 5510) && (pixel_index2 <= 5511)) || pixel_index2 == 5514 || ((pixel_index2 >= 5517) && (pixel_index2 <= 5520)) || ((pixel_index2 >= 5524) && (pixel_index2 <= 5532)) || ((pixel_index2 >= 5535) && (pixel_index2 <= 5537)) || ((pixel_index2 >= 5540) && (pixel_index2 <= 5541)) || pixel_index2 == 5544 || ((pixel_index2 >= 5548) && (pixel_index2 <= 5549)) || ((pixel_index2 >= 5553) && (pixel_index2 <= 5556)) || ((pixel_index2 >= 5560) && (pixel_index2 <= 5565)) || ((pixel_index2 >= 5570) && (pixel_index2 <= 5575)) || pixel_index2 == 5584 || pixel_index2 == 5587 || ((pixel_index2 >= 5590) && (pixel_index2 <= 5593)) || pixel_index2 == 5596 || pixel_index2 == 5603 || pixel_index2 == 5610 || pixel_index2 == 5613 || ((pixel_index2 >= 5620) && (pixel_index2 <= 5624)) || pixel_index2 == 5633 || pixel_index2 == 5640 || pixel_index2 == 5649 || ((pixel_index2 >= 5656) && (pixel_index2 <= 5661)) || ((pixel_index2 >= 5667) && (pixel_index2 <= 5671)) || pixel_index2 == 5680 || pixel_index2 == 5683 || ((pixel_index2 >= 5686) && (pixel_index2 <= 5689)) || pixel_index2 == 5692 || pixel_index2 == 5699 || pixel_index2 == 5706 || pixel_index2 == 5709 || ((pixel_index2 >= 5716) && (pixel_index2 <= 5720)) || pixel_index2 == 5729 || pixel_index2 == 5736 || pixel_index2 == 5745 || ((pixel_index2 >= 5752) && (pixel_index2 <= 5756)) || ((pixel_index2 >= 5763) && (pixel_index2 <= 5768)) || ((pixel_index2 >= 5775) && (pixel_index2 <= 5776)) || ((pixel_index2 >= 5778) && (pixel_index2 <= 5780)) || ((pixel_index2 >= 5782) && (pixel_index2 <= 5785)) || ((pixel_index2 >= 5787) && (pixel_index2 <= 5789)) || ((pixel_index2 >= 5794) && (pixel_index2 <= 5796)) || ((pixel_index2 >= 5801) && (pixel_index2 <= 5802)) || ((pixel_index2 >= 5804) && (pixel_index2 <= 5806)) || ((pixel_index2 >= 5811) && (pixel_index2 <= 5817)) || ((pixel_index2 >= 5824) && (pixel_index2 <= 5826)) || ((pixel_index2 >= 5831) && (pixel_index2 <= 5833)) || ((pixel_index2 >= 5840) && (pixel_index2 <= 5842)) || ((pixel_index2 >= 5847) && (pixel_index2 <= 5852)) || (pixel_index2 >= 5868) && (pixel_index2 <= 5940)) oled_data2 = 16'b0000000000001010;
                    else if (pixel_index2 == 323 || pixel_index2 == 327 || pixel_index2 == 331 || pixel_index2 == 335 || pixel_index2 == 339 || pixel_index2 == 419 || pixel_index2 == 423 || pixel_index2 == 427 || pixel_index2 == 431 || pixel_index2 == 435 || pixel_index2 == 3253 || pixel_index2 == 3349) oled_data2 = 16'b0000010100000000;
                    else if (pixel_index2 == 511 || pixel_index2 == 535 || pixel_index2 == 539 || pixel_index2 == 543 || pixel_index2 == 547 || pixel_index2 == 551 || pixel_index2 == 555 || pixel_index2 == 559 || pixel_index2 == 563 || pixel_index2 == 567 || pixel_index2 == 571 || pixel_index2 == 607 || pixel_index2 == 631 || pixel_index2 == 635 || pixel_index2 == 639 || pixel_index2 == 643 || pixel_index2 == 647 || pixel_index2 == 651 || pixel_index2 == 655 || pixel_index2 == 659 || pixel_index2 == 663 || pixel_index2 == 667 || pixel_index2 == 3488) oled_data2 = 16'b1010000000000000;
                    else if (pixel_index2 == 1086 || pixel_index2 == 1110 || pixel_index2 == 1114 || pixel_index2 == 1118 || pixel_index2 == 1122 || pixel_index2 == 1126 || pixel_index2 == 1130 || pixel_index2 == 1134 || pixel_index2 == 1138 || pixel_index2 == 1142 || pixel_index2 == 1146) oled_data2 = 16'b0000001010000000;
                    else if (pixel_index2 == 1090 || pixel_index2 == 1094 || pixel_index2 == 1098 || pixel_index2 == 1102 || pixel_index2 == 1106) oled_data2 = 16'b1111011110001010;
                    else if (((pixel_index2 >= 1281) && (pixel_index2 <= 1282)) || pixel_index2 == 1292 || pixel_index2 == 1295 || ((pixel_index2 >= 1297) && (pixel_index2 <= 1299)) || pixel_index2 == 1302 || ((pixel_index2 >= 1304) && (pixel_index2 <= 1305)) || pixel_index2 == 1307 || pixel_index2 == 1309 || pixel_index2 == 1311 || pixel_index2 == 1313 || pixel_index2 == 1377 || ((pixel_index2 >= 1392) && (pixel_index2 <= 1395)) || ((pixel_index2 >= 1397) && (pixel_index2 <= 1399)) || pixel_index2 == 1401 || ((pixel_index2 >= 1403) && (pixel_index2 <= 1404)) || pixel_index2 == 1406 || pixel_index2 == 1409 || ((pixel_index2 >= 1487) && (pixel_index2 <= 1488)) || pixel_index2 == 1490 || pixel_index2 == 1493 || pixel_index2 == 1495 || pixel_index2 == 1497 || ((pixel_index2 >= 1499) && (pixel_index2 <= 1500)) || ((pixel_index2 >= 1502) && (pixel_index2 <= 1503)) || pixel_index2 == 1505 || pixel_index2 == 1697 || pixel_index2 == 1776 || ((pixel_index2 >= 1790) && (pixel_index2 <= 1791)) || pixel_index2 == 1793 || pixel_index2 == 1817 || pixel_index2 == 1871 || pixel_index2 == 1914 || pixel_index2 == 1974 || ((pixel_index2 >= 1989) && (pixel_index2 <= 1990)) || pixel_index2 == 1992 || pixel_index2 == 1995 || ((pixel_index2 >= 1997) && (pixel_index2 <= 1999)) || ((pixel_index2 >= 2009) && (pixel_index2 <= 2010)) || pixel_index2 == 2047 || ((pixel_index2 >= 2070) && (pixel_index2 <= 2071)) || pixel_index2 == 2083 || ((pixel_index2 >= 2086) && (pixel_index2 <= 2088)) || pixel_index2 == 2090 || pixel_index2 == 2094 || pixel_index2 == 2106 || pixel_index2 == 2141 || pixel_index2 == 2143 || ((pixel_index2 >= 2155) && (pixel_index2 <= 2156)) || pixel_index2 == 2179 || ((pixel_index2 >= 2185) && (pixel_index2 <= 2187)) || pixel_index2 == 2189 || pixel_index2 == 2240 || pixel_index2 == 2243 || pixel_index2 == 2251 || pixel_index2 == 2336 || pixel_index2 == 2338 || pixel_index2 == 2340 || pixel_index2 == 2548 || ((pixel_index2 >= 2550) && (pixel_index2 <= 2551)) || ((pixel_index2 >= 2562) && (pixel_index2 <= 2563)) || ((pixel_index2 >= 2567) && (pixel_index2 <= 2579)) || ((pixel_index2 >= 2645) && (pixel_index2 <= 2646)) || pixel_index2 == 2658 || pixel_index2 == 2660 || ((pixel_index2 >= 2663) && (pixel_index2 <= 2675)) || ((pixel_index2 >= 2759) && (pixel_index2 <= 2771)) || ((pixel_index2 >= 2925) && (pixel_index2 <= 2926)) || pixel_index2 == 2937 || pixel_index2 == 2946 || pixel_index2 == 3022 || ((pixel_index2 >= 3105) && (pixel_index2 <= 3106)) || pixel_index2 == 3201 || pixel_index2 == 3217 || ((pixel_index2 >= 3230) && (pixel_index2 <= 3231)) || pixel_index2 == 3313 || pixel_index2 == 3324 || pixel_index2 == 3408 || ((pixel_index2 >= 3421) && (pixel_index2 <= 3422)) || ((pixel_index2 >= 3503) && (pixel_index2 <= 3504)) || ((pixel_index2 >= 3533) && (pixel_index2 <= 3536)) || pixel_index2 == 3629 || pixel_index2 == 3632) oled_data2 = 16'b1010010100010100;
                    else if (pixel_index2 == 1287 || pixel_index2 == 1289 || pixel_index2 == 1479 || pixel_index2 == 1481 || pixel_index2 == 1667 || pixel_index2 == 1669 || pixel_index2 == 1671 || pixel_index2 == 1673 || pixel_index2 == 1675 || pixel_index2 == 1677 || pixel_index2 == 1859 || pixel_index2 == 1861 || pixel_index2 == 1863 || pixel_index2 == 1865 || pixel_index2 == 1867 || pixel_index2 == 1869 || ((pixel_index2 >= 1879) && (pixel_index2 <= 1881)) || ((pixel_index2 >= 1889) && (pixel_index2 <= 1891)) || ((pixel_index2 >= 1975) && (pixel_index2 <= 1987)) || ((pixel_index2 >= 2002) && (pixel_index2 <= 2007)) || pixel_index2 == 2055 || pixel_index2 == 2057 || ((pixel_index2 >= 2072) && (pixel_index2 <= 2073)) || ((pixel_index2 >= 2081) && (pixel_index2 <= 2082)) || ((pixel_index2 >= 2097) && (pixel_index2 <= 2103)) || pixel_index2 == 2169 || pixel_index2 == 2177 || ((pixel_index2 >= 2193) && (pixel_index2 <= 2194)) || ((pixel_index2 >= 2198) && (pixel_index2 <= 2199)) || pixel_index2 == 2239 || ((pixel_index2 >= 2241) && (pixel_index2 <= 2242)) || pixel_index2 == 2244 || pixel_index2 == 2247 || pixel_index2 == 2249 || pixel_index2 == 2265 || pixel_index2 == 2273 || ((pixel_index2 >= 2289) && (pixel_index2 <= 2290)) || ((pixel_index2 >= 2294) && (pixel_index2 <= 2295)) || pixel_index2 == 2335 || pixel_index2 == 2337 || pixel_index2 == 2339 || ((pixel_index2 >= 2356) && (pixel_index2 <= 2361)) || ((pixel_index2 >= 2369) && (pixel_index2 <= 2373)) || ((pixel_index2 >= 2385) && (pixel_index2 <= 2391)) || ((pixel_index2 >= 2438) && (pixel_index2 <= 2442)) || ((pixel_index2 >= 2452) && (pixel_index2 <= 2457)) || ((pixel_index2 >= 2465) && (pixel_index2 <= 2469)) || ((pixel_index2 >= 2481) && (pixel_index2 <= 2486)) || pixel_index2 == 2533 || pixel_index2 == 2539 || pixel_index2 == 2549 || ((pixel_index2 >= 2552) && (pixel_index2 <= 2553)) || pixel_index2 == 2561 || ((pixel_index2 >= 2564) && (pixel_index2 <= 2565)) || ((pixel_index2 >= 2627) && (pixel_index2 <= 2629)) || pixel_index2 == 2635 || ((pixel_index2 >= 2637) && (pixel_index2 <= 2638)) || pixel_index2 == 2649 || pixel_index2 == 2657 || ((pixel_index2 >= 2722) && (pixel_index2 <= 2725)) || pixel_index2 == 2731 || ((pixel_index2 >= 2733) && (pixel_index2 <= 2734)) || ((pixel_index2 >= 2743) && (pixel_index2 <= 2755)) || ((pixel_index2 >= 2818) && (pixel_index2 <= 2821)) || pixel_index2 == 2827 || ((pixel_index2 >= 2829) && (pixel_index2 <= 2830)) || ((pixel_index2 >= 2839) && (pixel_index2 <= 2841)) || ((pixel_index2 >= 2849) && (pixel_index2 <= 2851)) || ((pixel_index2 >= 2914) && (pixel_index2 <= 2917)) || pixel_index2 == 2923 || pixel_index2 == 2936 || pixel_index2 == 2945 || pixel_index2 == 2963 || ((pixel_index2 >= 3014) && (pixel_index2 <= 3018)) || ((pixel_index2 >= 3061) && (pixel_index2 <= 3062)) || pixel_index2 == 3064 || ((pixel_index2 >= 3108) && (pixel_index2 <= 3116)) || pixel_index2 == 3160 || ((pixel_index2 >= 3204) && (pixel_index2 <= 3212)) || ((pixel_index2 >= 3300) && (pixel_index2 <= 3308)) || pixel_index2 == 3317 || ((pixel_index2 >= 3319) && (pixel_index2 <= 3320)) || ((pixel_index2 >= 3330) && (pixel_index2 <= 3331)) || pixel_index2 == 3333 || pixel_index2 == 3338 || ((pixel_index2 >= 3396) && (pixel_index2 <= 3404)) || pixel_index2 == 3433 || ((pixel_index2 >= 3436) && (pixel_index2 <= 3437)) || ((pixel_index2 >= 3492) && (pixel_index2 <= 3500)) || ((pixel_index2 >= 3588) && (pixel_index2 <= 3596)) || ((pixel_index2 >= 3684) && (pixel_index2 <= 3692)) || ((pixel_index2 >= 3724) && (pixel_index2 <= 3729)) || ((pixel_index2 >= 3820) && (pixel_index2 <= 3825)) || ((pixel_index2 >= 3893) && (pixel_index2 <= 3894)) || ((pixel_index2 >= 3897) && (pixel_index2 <= 3905)) || ((pixel_index2 >= 3908) && (pixel_index2 <= 3909)) || ((pixel_index2 >= 3989) && (pixel_index2 <= 3990)) || ((pixel_index2 >= 3994) && (pixel_index2 <= 4000)) || ((pixel_index2 >= 4004) && (pixel_index2 <= 4005)) || ((pixel_index2 >= 4085) && (pixel_index2 <= 4086)) || ((pixel_index2 >= 4090) && (pixel_index2 <= 4096)) || ((pixel_index2 >= 4100) && (pixel_index2 <= 4101)) || pixel_index2 == 4706 || pixel_index2 == 4797 || pixel_index2 == 5666 || pixel_index2 == 5757) oled_data2 = 16'b0101001010001010;
                    else if (pixel_index2 == 1296 || ((pixel_index2 >= 1300) && (pixel_index2 <= 1301)) || pixel_index2 == 1303 || pixel_index2 == 1306 || pixel_index2 == 1308 || pixel_index2 == 1310 || pixel_index2 == 1312 || pixel_index2 == 1391 || pixel_index2 == 1396 || pixel_index2 == 1400 || pixel_index2 == 1402 || pixel_index2 == 1405 || ((pixel_index2 >= 1407) && (pixel_index2 <= 1408)) || pixel_index2 == 1489 || ((pixel_index2 >= 1491) && (pixel_index2 <= 1492)) || pixel_index2 == 1494 || pixel_index2 == 1496 || pixel_index2 == 1498 || pixel_index2 == 1501 || pixel_index2 == 1504 || pixel_index2 == 3353 || pixel_index2 == 3449 || pixel_index2 == 3545) oled_data2 = 16'b0101001010010100;
                    else if (((pixel_index2 >= 1317) && (pixel_index2 <= 1319)) || pixel_index2 == 1322 || pixel_index2 == 1324 || pixel_index2 == 1327 || pixel_index2 == 1329 || pixel_index2 == 1332 || pixel_index2 == 1334 || pixel_index2 == 1415 || pixel_index2 == 1418 || pixel_index2 == 1420 || pixel_index2 == 1423 || pixel_index2 == 1425 || pixel_index2 == 1428 || pixel_index2 == 1430 || pixel_index2 == 1511 || ((pixel_index2 >= 1514) && (pixel_index2 <= 1516)) || ((pixel_index2 >= 1519) && (pixel_index2 <= 1521)) || pixel_index2 == 1607 || pixel_index2 == 1615 || pixel_index2 == 1617 || pixel_index2 == 1703 || ((pixel_index2 >= 1711) && (pixel_index2 <= 1713)) || (pixel_index2 >= 1716) && (pixel_index2 <= 1718)) oled_data2 = 16'b1010000000001010;
                    else if (((pixel_index2 >= 1574) && (pixel_index2 <= 1578)) || pixel_index2 == 1670 || pixel_index2 == 1674 || pixel_index2 == 1766 || pixel_index2 == 1770 || pixel_index2 == 1862 || pixel_index2 == 1866 || ((pixel_index2 >= 1958) && (pixel_index2 <= 1962)) || ((pixel_index2 >= 3938) && (pixel_index2 <= 3939)) || pixel_index2 == 3942 || pixel_index2 == 3945 || ((pixel_index2 >= 3947) && (pixel_index2 <= 3950)) || pixel_index2 == 3952 || ((pixel_index2 >= 3954) && (pixel_index2 <= 3955)) || ((pixel_index2 >= 3959) && (pixel_index2 <= 3962)) || ((pixel_index2 >= 3964) && (pixel_index2 <= 3967)) || ((pixel_index2 >= 3969) && (pixel_index2 <= 3972)) || ((pixel_index2 >= 3974) && (pixel_index2 <= 3977)) || pixel_index2 == 3979 || ((pixel_index2 >= 3981) && (pixel_index2 <= 3982)) || ((pixel_index2 >= 3984) && (pixel_index2 <= 3986)) || ((pixel_index2 >= 4034) && (pixel_index2 <= 4035)) || ((pixel_index2 >= 4039) && (pixel_index2 <= 4040)) || ((pixel_index2 >= 4045) && (pixel_index2 <= 4046)) || pixel_index2 == 4048 || ((pixel_index2 >= 4050) && (pixel_index2 <= 4051)) || ((pixel_index2 >= 4057) && (pixel_index2 <= 4058)) || ((pixel_index2 >= 4060) && (pixel_index2 <= 4061)) || pixel_index2 == 4065 || ((pixel_index2 >= 4067) && (pixel_index2 <= 4068)) || pixel_index2 == 4070 || ((pixel_index2 >= 4072) && (pixel_index2 <= 4073)) || ((pixel_index2 >= 4075) && (pixel_index2 <= 4078)) || ((pixel_index2 >= 4082) && (pixel_index2 <= 4083)) || ((pixel_index2 >= 4130) && (pixel_index2 <= 4131)) || ((pixel_index2 >= 4135) && (pixel_index2 <= 4136)) || ((pixel_index2 >= 4139) && (pixel_index2 <= 4140)) || pixel_index2 == 4142 || pixel_index2 == 4144 || ((pixel_index2 >= 4146) && (pixel_index2 <= 4147)) || ((pixel_index2 >= 4151) && (pixel_index2 <= 4152)) || pixel_index2 == 4154 || ((pixel_index2 >= 4157) && (pixel_index2 <= 4159)) || pixel_index2 == 4161 || ((pixel_index2 >= 4163) && (pixel_index2 <= 4164)) || pixel_index2 == 4166 || ((pixel_index2 >= 4168) && (pixel_index2 <= 4169)) || pixel_index2 == 4171 || ((pixel_index2 >= 4173) && (pixel_index2 <= 4174)) || ((pixel_index2 >= 4178) && (pixel_index2 <= 4179)) || ((pixel_index2 >= 4225) && (pixel_index2 <= 4228)) || pixel_index2 == 4230 || pixel_index2 == 4233 || ((pixel_index2 >= 4235) && (pixel_index2 <= 4238)) || ((pixel_index2 >= 4240) && (pixel_index2 <= 4243)) || ((pixel_index2 >= 4247) && (pixel_index2 <= 4250)) || ((pixel_index2 >= 4252) && (pixel_index2 <= 4254)) || ((pixel_index2 >= 4257) && (pixel_index2 <= 4260)) || ((pixel_index2 >= 4262) && (pixel_index2 <= 4265)) || pixel_index2 == 4267 || ((pixel_index2 >= 4269) && (pixel_index2 <= 4270)) || (pixel_index2 >= 4272) && (pixel_index2 <= 4274)) oled_data2 = 16'b1111001010010100;
                    else if (pixel_index2 == 3229 || (pixel_index2 >= 3325) && (pixel_index2 <= 3326)) oled_data2 = 16'b0101010100001010;
                    else if (pixel_index2 == 3394 || pixel_index2 == 3490) oled_data2 = 16'b0000000000010100;
                    else if (pixel_index2 == 3532 || pixel_index2 == 3537) oled_data2 = 16'b0101000000000000;
                    else if (((pixel_index2 >= 4423) && (pixel_index2 <= 4505)) || ((pixel_index2 >= 4513) && (pixel_index2 <= 4518)) || (pixel_index2 >= 4602) && (pixel_index2 <= 4606)) oled_data2 = 16'b0000001010011110;
                    else if (((pixel_index2 >= 4519) && (pixel_index2 <= 4601)) || ((pixel_index2 >= 4609) && (pixel_index2 <= 4619)) || ((pixel_index2 >= 4693) && (pixel_index2 <= 4702)) || pixel_index2 == 4705 || pixel_index2 == 4798 || pixel_index2 == 4801 || pixel_index2 == 4894 || ((pixel_index2 >= 4897) && (pixel_index2 <= 4898)) || ((pixel_index2 >= 4989) && (pixel_index2 <= 4990)) || pixel_index2 == 4993 || pixel_index2 == 5086 || pixel_index2 == 5089 || pixel_index2 == 5182 || pixel_index2 == 5185 || pixel_index2 == 5278 || pixel_index2 == 5281 || pixel_index2 == 5374 || pixel_index2 == 5377 || pixel_index2 == 5470 || pixel_index2 == 5473 || pixel_index2 == 5566 || pixel_index2 == 5569 || pixel_index2 == 5662 || pixel_index2 == 5665 || pixel_index2 == 5758 || pixel_index2 == 5761 || pixel_index2 == 5854 || ((pixel_index2 >= 5857) && (pixel_index2 <= 5867)) || ((pixel_index2 >= 5941) && (pixel_index2 <= 5950)) || (pixel_index2 >= 5959) && (pixel_index2 <= 6041)) oled_data2 = 16'b0000001010010100;
                    else if (pixel_index2 == 4813 || pixel_index2 == 4818 || ((pixel_index2 >= 4821) && (pixel_index2 <= 4826)) || ((pixel_index2 >= 4830) && (pixel_index2 <= 4833)) || ((pixel_index2 >= 4836) && (pixel_index2 <= 4837)) || pixel_index2 == 4840 || pixel_index2 == 4844 || ((pixel_index2 >= 4847) && (pixel_index2 <= 4850)) || pixel_index2 == 4862 || ((pixel_index2 >= 4866) && (pixel_index2 <= 4867)) || pixel_index2 == 4870 || ((pixel_index2 >= 4874) && (pixel_index2 <= 4879)) || ((pixel_index2 >= 4883) && (pixel_index2 <= 4886)) || pixel_index2 == 4908 || pixel_index2 == 4913 || pixel_index2 == 4916 || pixel_index2 == 4923 || pixel_index2 == 4925 || pixel_index2 == 4930 || pixel_index2 == 4934 || pixel_index2 == 4937 || pixel_index2 == 4939 || pixel_index2 == 4942 || pixel_index2 == 4947 || pixel_index2 == 4957 || pixel_index2 == 4964 || pixel_index2 == 4967 || pixel_index2 == 4969 || pixel_index2 == 4976 || pixel_index2 == 4978 || pixel_index2 == 4983 || pixel_index2 == 5031 || pixel_index2 == 5061 || pixel_index2 == 5221 || pixel_index2 == 5251 || ((pixel_index2 >= 5268) && (pixel_index2 <= 5270)) || pixel_index2 == 5316 || pixel_index2 == 5346 || pixel_index2 == 5367 || pixel_index2 == 5504 || pixel_index2 == 5521 || pixel_index2 == 5547 || pixel_index2 == 5550 || pixel_index2 == 5557 || ((pixel_index2 >= 5576) && (pixel_index2 <= 5579)) || ((pixel_index2 >= 5582) && (pixel_index2 <= 5583)) || ((pixel_index2 >= 5597) && (pixel_index2 <= 5599)) || ((pixel_index2 >= 5606) && (pixel_index2 <= 5607)) || ((pixel_index2 >= 5614) && (pixel_index2 <= 5616)) || ((pixel_index2 >= 5625) && (pixel_index2 <= 5628)) || ((pixel_index2 >= 5631) && (pixel_index2 <= 5632)) || ((pixel_index2 >= 5636) && (pixel_index2 <= 5637)) || ((pixel_index2 >= 5644) && (pixel_index2 <= 5645)) || (pixel_index2 >= 5650) && (pixel_index2 <= 5652)) oled_data2 = 16'b0101001010000000;
                    else if (pixel_index2 == 4909 || pixel_index2 == 4914 || ((pixel_index2 >= 4917) && (pixel_index2 <= 4922)) || ((pixel_index2 >= 4926) && (pixel_index2 <= 4929)) || ((pixel_index2 >= 4932) && (pixel_index2 <= 4933)) || pixel_index2 == 4936 || pixel_index2 == 4940 || ((pixel_index2 >= 4943) && (pixel_index2 <= 4946)) || pixel_index2 == 4958 || ((pixel_index2 >= 4962) && (pixel_index2 <= 4963)) || pixel_index2 == 4966 || ((pixel_index2 >= 4970) && (pixel_index2 <= 4975)) || ((pixel_index2 >= 4979) && (pixel_index2 <= 4982)) || ((pixel_index2 >= 5004) && (pixel_index2 <= 5005)) || ((pixel_index2 >= 5009) && (pixel_index2 <= 5010)) || ((pixel_index2 >= 5012) && (pixel_index2 <= 5019)) || ((pixel_index2 >= 5021) && (pixel_index2 <= 5026)) || ((pixel_index2 >= 5028) && (pixel_index2 <= 5030)) || ((pixel_index2 >= 5032) && (pixel_index2 <= 5033)) || ((pixel_index2 >= 5035) && (pixel_index2 <= 5036)) || ((pixel_index2 >= 5038) && (pixel_index2 <= 5043)) || ((pixel_index2 >= 5053) && (pixel_index2 <= 5054)) || ((pixel_index2 >= 5058) && (pixel_index2 <= 5060)) || ((pixel_index2 >= 5062) && (pixel_index2 <= 5063)) || ((pixel_index2 >= 5065) && (pixel_index2 <= 5072)) || ((pixel_index2 >= 5074) && (pixel_index2 <= 5079)) || ((pixel_index2 >= 5100) && (pixel_index2 <= 5101)) || ((pixel_index2 >= 5105) && (pixel_index2 <= 5106)) || ((pixel_index2 >= 5108) && (pixel_index2 <= 5110)) || ((pixel_index2 >= 5113) && (pixel_index2 <= 5115)) || ((pixel_index2 >= 5120) && (pixel_index2 <= 5122)) || ((pixel_index2 >= 5125) && (pixel_index2 <= 5129)) || ((pixel_index2 >= 5131) && (pixel_index2 <= 5132)) || ((pixel_index2 >= 5137) && (pixel_index2 <= 5139)) || ((pixel_index2 >= 5149) && (pixel_index2 <= 5150)) || ((pixel_index2 >= 5155) && (pixel_index2 <= 5159)) || ((pixel_index2 >= 5161) && (pixel_index2 <= 5163)) || ((pixel_index2 >= 5166) && (pixel_index2 <= 5168)) || ((pixel_index2 >= 5170) && (pixel_index2 <= 5172)) || ((pixel_index2 >= 5196) && (pixel_index2 <= 5197)) || ((pixel_index2 >= 5201) && (pixel_index2 <= 5202)) || ((pixel_index2 >= 5204) && (pixel_index2 <= 5205)) || ((pixel_index2 >= 5210) && (pixel_index2 <= 5211)) || ((pixel_index2 >= 5217) && (pixel_index2 <= 5218)) || ((pixel_index2 >= 5222) && (pixel_index2 <= 5225)) || ((pixel_index2 >= 5227) && (pixel_index2 <= 5228)) || ((pixel_index2 >= 5234) && (pixel_index2 <= 5235)) || ((pixel_index2 >= 5245) && (pixel_index2 <= 5246)) || ((pixel_index2 >= 5252) && (pixel_index2 <= 5255)) || ((pixel_index2 >= 5257) && (pixel_index2 <= 5258)) || ((pixel_index2 >= 5263) && (pixel_index2 <= 5264)) || ((pixel_index2 >= 5266) && (pixel_index2 <= 5267)) || ((pixel_index2 >= 5292) && (pixel_index2 <= 5293)) || ((pixel_index2 >= 5297) && (pixel_index2 <= 5298)) || ((pixel_index2 >= 5300) && (pixel_index2 <= 5301)) || ((pixel_index2 >= 5306) && (pixel_index2 <= 5307)) || ((pixel_index2 >= 5313) && (pixel_index2 <= 5314)) || ((pixel_index2 >= 5317) && (pixel_index2 <= 5321)) || ((pixel_index2 >= 5323) && (pixel_index2 <= 5324)) || ((pixel_index2 >= 5330) && (pixel_index2 <= 5331)) || ((pixel_index2 >= 5341) && (pixel_index2 <= 5342)) || ((pixel_index2 >= 5347) && (pixel_index2 <= 5351)) || ((pixel_index2 >= 5353) && (pixel_index2 <= 5354)) || ((pixel_index2 >= 5359) && (pixel_index2 <= 5360)) || ((pixel_index2 >= 5362) && (pixel_index2 <= 5366)) || ((pixel_index2 >= 5388) && (pixel_index2 <= 5389)) || ((pixel_index2 >= 5393) && (pixel_index2 <= 5394)) || ((pixel_index2 >= 5396) && (pixel_index2 <= 5397)) || ((pixel_index2 >= 5402) && (pixel_index2 <= 5403)) || ((pixel_index2 >= 5409) && (pixel_index2 <= 5410)) || ((pixel_index2 >= 5412) && (pixel_index2 <= 5414)) || ((pixel_index2 >= 5416) && (pixel_index2 <= 5417)) || ((pixel_index2 >= 5419) && (pixel_index2 <= 5420)) || ((pixel_index2 >= 5426) && (pixel_index2 <= 5427)) || ((pixel_index2 >= 5437) && (pixel_index2 <= 5438)) || ((pixel_index2 >= 5442) && (pixel_index2 <= 5444)) || ((pixel_index2 >= 5446) && (pixel_index2 <= 5447)) || ((pixel_index2 >= 5449) && (pixel_index2 <= 5450)) || ((pixel_index2 >= 5455) && (pixel_index2 <= 5456)) || ((pixel_index2 >= 5459) && (pixel_index2 <= 5463)) || ((pixel_index2 >= 5484) && (pixel_index2 <= 5485)) || ((pixel_index2 >= 5489) && (pixel_index2 <= 5490)) || ((pixel_index2 >= 5492) && (pixel_index2 <= 5493)) || ((pixel_index2 >= 5498) && (pixel_index2 <= 5499)) || ((pixel_index2 >= 5505) && (pixel_index2 <= 5506)) || ((pixel_index2 >= 5508) && (pixel_index2 <= 5509)) || ((pixel_index2 >= 5512) && (pixel_index2 <= 5513)) || ((pixel_index2 >= 5515) && (pixel_index2 <= 5516)) || ((pixel_index2 >= 5522) && (pixel_index2 <= 5523)) || ((pixel_index2 >= 5533) && (pixel_index2 <= 5534)) || ((pixel_index2 >= 5538) && (pixel_index2 <= 5539)) || ((pixel_index2 >= 5542) && (pixel_index2 <= 5543)) || ((pixel_index2 >= 5545) && (pixel_index2 <= 5546)) || ((pixel_index2 >= 5551) && (pixel_index2 <= 5552)) || ((pixel_index2 >= 5558) && (pixel_index2 <= 5559)) || ((pixel_index2 >= 5580) && (pixel_index2 <= 5581)) || ((pixel_index2 >= 5585) && (pixel_index2 <= 5586)) || ((pixel_index2 >= 5588) && (pixel_index2 <= 5589)) || ((pixel_index2 >= 5594) && (pixel_index2 <= 5595)) || ((pixel_index2 >= 5600) && (pixel_index2 <= 5602)) || ((pixel_index2 >= 5604) && (pixel_index2 <= 5605)) || ((pixel_index2 >= 5608) && (pixel_index2 <= 5609)) || ((pixel_index2 >= 5611) && (pixel_index2 <= 5612)) || ((pixel_index2 >= 5617) && (pixel_index2 <= 5619)) || ((pixel_index2 >= 5629) && (pixel_index2 <= 5630)) || ((pixel_index2 >= 5634) && (pixel_index2 <= 5635)) || ((pixel_index2 >= 5638) && (pixel_index2 <= 5639)) || ((pixel_index2 >= 5641) && (pixel_index2 <= 5643)) || ((pixel_index2 >= 5646) && (pixel_index2 <= 5648)) || ((pixel_index2 >= 5653) && (pixel_index2 <= 5655)) || ((pixel_index2 >= 5672) && (pixel_index2 <= 5679)) || ((pixel_index2 >= 5681) && (pixel_index2 <= 5682)) || ((pixel_index2 >= 5684) && (pixel_index2 <= 5685)) || ((pixel_index2 >= 5690) && (pixel_index2 <= 5691)) || ((pixel_index2 >= 5693) && (pixel_index2 <= 5698)) || ((pixel_index2 >= 5700) && (pixel_index2 <= 5705)) || ((pixel_index2 >= 5707) && (pixel_index2 <= 5708)) || ((pixel_index2 >= 5710) && (pixel_index2 <= 5715)) || ((pixel_index2 >= 5721) && (pixel_index2 <= 5728)) || ((pixel_index2 >= 5730) && (pixel_index2 <= 5735)) || ((pixel_index2 >= 5737) && (pixel_index2 <= 5744)) || ((pixel_index2 >= 5746) && (pixel_index2 <= 5751)) || ((pixel_index2 >= 5769) && (pixel_index2 <= 5774)) || pixel_index2 == 5777 || pixel_index2 == 5781 || pixel_index2 == 5786 || ((pixel_index2 >= 5790) && (pixel_index2 <= 5793)) || ((pixel_index2 >= 5797) && (pixel_index2 <= 5800)) || pixel_index2 == 5803 || ((pixel_index2 >= 5807) && (pixel_index2 <= 5810)) || ((pixel_index2 >= 5818) && (pixel_index2 <= 5823)) || ((pixel_index2 >= 5827) && (pixel_index2 <= 5830)) || ((pixel_index2 >= 5834) && (pixel_index2 <= 5839)) || (pixel_index2 >= 5843) && (pixel_index2 <= 5846)) oled_data2 = 16'b1111010100010100;
                    else oled_data2 = 0;
                end
                3: begin
                    if (pixel_index2 == 97 || pixel_index2 == 99 || pixel_index2 == 101 || ((pixel_index2 >= 103) && (pixel_index2 <= 104)) || ((pixel_index2 >= 106) && (pixel_index2 <= 109)) || pixel_index2 == 111 || ((pixel_index2 >= 113) && (pixel_index2 <= 114)) || ((pixel_index2 >= 118) && (pixel_index2 <= 120)) || pixel_index2 == 195 || pixel_index2 == 197 || ((pixel_index2 >= 199) && (pixel_index2 <= 200)) || pixel_index2 == 202 || ((pixel_index2 >= 204) && (pixel_index2 <= 205)) || pixel_index2 == 207 || ((pixel_index2 >= 209) && (pixel_index2 <= 210)) || pixel_index2 == 213 || pixel_index2 == 289 || ((pixel_index2 >= 291) && (pixel_index2 <= 296)) || pixel_index2 == 298 || ((pixel_index2 >= 300) && (pixel_index2 <= 301)) || pixel_index2 == 303 || ((pixel_index2 >= 305) && (pixel_index2 <= 306)) || ((pixel_index2 >= 310) && (pixel_index2 <= 312)) || pixel_index2 == 385 || ((pixel_index2 >= 387) && (pixel_index2 <= 392)) || pixel_index2 == 394 || ((pixel_index2 >= 396) && (pixel_index2 <= 397)) || ((pixel_index2 >= 399) && (pixel_index2 <= 402)) || pixel_index2 == 408 || ((pixel_index2 >= 501) && (pixel_index2 <= 504)) || ((pixel_index2 >= 674) && (pixel_index2 <= 675)) || ((pixel_index2 >= 678) && (pixel_index2 <= 681)) || ((pixel_index2 >= 685) && (pixel_index2 <= 686)) || pixel_index2 == 688 || ((pixel_index2 >= 690) && (pixel_index2 <= 691)) || ((pixel_index2 >= 693) && (pixel_index2 <= 696)) || ((pixel_index2 >= 770) && (pixel_index2 <= 771)) || pixel_index2 == 774 || ((pixel_index2 >= 776) && (pixel_index2 <= 777)) || ((pixel_index2 >= 779) && (pixel_index2 <= 782)) || pixel_index2 == 784 || ((pixel_index2 >= 786) && (pixel_index2 <= 787)) || ((pixel_index2 >= 790) && (pixel_index2 <= 791)) || ((pixel_index2 >= 866) && (pixel_index2 <= 867)) || pixel_index2 == 870 || ((pixel_index2 >= 872) && (pixel_index2 <= 873)) || pixel_index2 == 875 || ((pixel_index2 >= 877) && (pixel_index2 <= 878)) || pixel_index2 == 880 || ((pixel_index2 >= 882) && (pixel_index2 <= 883)) || ((pixel_index2 >= 886) && (pixel_index2 <= 887)) || ((pixel_index2 >= 895) && (pixel_index2 <= 896)) || ((pixel_index2 >= 899) && (pixel_index2 <= 900)) || ((pixel_index2 >= 903) && (pixel_index2 <= 904)) || ((pixel_index2 >= 907) && (pixel_index2 <= 908)) || ((pixel_index2 >= 911) && (pixel_index2 <= 912)) || ((pixel_index2 >= 915) && (pixel_index2 <= 916)) || ((pixel_index2 >= 919) && (pixel_index2 <= 920)) || ((pixel_index2 >= 923) && (pixel_index2 <= 924)) || ((pixel_index2 >= 927) && (pixel_index2 <= 928)) || ((pixel_index2 >= 931) && (pixel_index2 <= 932)) || ((pixel_index2 >= 935) && (pixel_index2 <= 936)) || ((pixel_index2 >= 939) && (pixel_index2 <= 940)) || ((pixel_index2 >= 943) && (pixel_index2 <= 944)) || ((pixel_index2 >= 947) && (pixel_index2 <= 948)) || ((pixel_index2 >= 951) && (pixel_index2 <= 952)) || ((pixel_index2 >= 955) && (pixel_index2 <= 956)) || ((pixel_index2 >= 961) && (pixel_index2 <= 964)) || pixel_index2 == 966 || ((pixel_index2 >= 968) && (pixel_index2 <= 969)) || ((pixel_index2 >= 971) && (pixel_index2 <= 974)) || ((pixel_index2 >= 976) && (pixel_index2 <= 979)) || ((pixel_index2 >= 981) && (pixel_index2 <= 984)) || ((pixel_index2 >= 1637) && (pixel_index2 <= 1638)) || ((pixel_index2 >= 1641) && (pixel_index2 <= 1644)) || ((pixel_index2 >= 1646) && (pixel_index2 <= 1649)) || ((pixel_index2 >= 1652) && (pixel_index2 <= 1654)) || pixel_index2 == 1732 || pixel_index2 == 1735 || pixel_index2 == 1740 || pixel_index2 == 1745 || pixel_index2 == 1747 || pixel_index2 == 1831 || pixel_index2 == 1836 || ((pixel_index2 >= 1839) && (pixel_index2 <= 1841)) || ((pixel_index2 >= 1844) && (pixel_index2 <= 1845)) || pixel_index2 == 1924 || pixel_index2 == 1927 || pixel_index2 == 1932 || pixel_index2 == 1937 || pixel_index2 == 1942 || ((pixel_index2 >= 2021) && (pixel_index2 <= 2022)) || pixel_index2 == 2028 || ((pixel_index2 >= 2030) && (pixel_index2 <= 2033)) || ((pixel_index2 >= 2035) && (pixel_index2 <= 2037)) || pixel_index2 == 2213 || pixel_index2 == 2216 || ((pixel_index2 >= 2219) && (pixel_index2 <= 2221)) || pixel_index2 == 2223 || pixel_index2 == 2226 || ((pixel_index2 >= 2228) && (pixel_index2 <= 2230)) || pixel_index2 == 2310 || pixel_index2 == 2312 || pixel_index2 == 2314 || pixel_index2 == 2319 || pixel_index2 == 2322 || pixel_index2 == 2325 || ((pixel_index2 >= 2406) && (pixel_index2 <= 2408)) || ((pixel_index2 >= 2411) && (pixel_index2 <= 2412)) || ((pixel_index2 >= 2415) && (pixel_index2 <= 2416)) || pixel_index2 == 2418 || pixel_index2 == 2421 || pixel_index2 == 2501 || pixel_index2 == 2504 || pixel_index2 == 2509 || pixel_index2 == 2511 || ((pixel_index2 >= 2513) && (pixel_index2 <= 2514)) || pixel_index2 == 2517 || ((pixel_index2 >= 2598) && (pixel_index2 <= 2600)) || ((pixel_index2 >= 2602) && (pixel_index2 <= 2604)) || pixel_index2 == 2607 || pixel_index2 == 2610 || ((pixel_index2 >= 2612) && (pixel_index2 <= 2614)) || pixel_index2 == 2788 || pixel_index2 == 2791 || ((pixel_index2 >= 2794) && (pixel_index2 <= 2795)) || ((pixel_index2 >= 2799) && (pixel_index2 <= 2800)) || ((pixel_index2 >= 2804) && (pixel_index2 <= 2805)) || pixel_index2 == 2885 || pixel_index2 == 2887 || pixel_index2 == 2889 || pixel_index2 == 2892 || pixel_index2 == 2894 || pixel_index2 == 2897 || pixel_index2 == 2899 || pixel_index2 == 2902 || ((pixel_index2 >= 2982) && (pixel_index2 <= 2983)) || pixel_index2 == 2988 || pixel_index2 == 2990 || pixel_index2 == 2993 || pixel_index2 == 2998 || pixel_index2 == 3077 || pixel_index2 == 3079 || pixel_index2 == 3081 || pixel_index2 == 3084 || pixel_index2 == 3086 || pixel_index2 == 3089 || pixel_index2 == 3091 || pixel_index2 == 3094 || ((pixel_index2 >= 3133) && (pixel_index2 <= 3134)) || pixel_index2 == 3172 || pixel_index2 == 3175 || ((pixel_index2 >= 3178) && (pixel_index2 <= 3179)) || ((pixel_index2 >= 3183) && (pixel_index2 <= 3184)) || ((pixel_index2 >= 3188) && (pixel_index2 <= 3189)) || pixel_index2 == 3228 || pixel_index2 == 3327 || ((pixel_index2 >= 3630) && (pixel_index2 <= 3631)) || ((pixel_index2 >= 3938) && (pixel_index2 <= 3939)) || pixel_index2 == 3942 || pixel_index2 == 3945 || ((pixel_index2 >= 3947) && (pixel_index2 <= 3950)) || pixel_index2 == 3952 || ((pixel_index2 >= 3954) && (pixel_index2 <= 3955)) || ((pixel_index2 >= 3959) && (pixel_index2 <= 3962)) || ((pixel_index2 >= 3964) && (pixel_index2 <= 3967)) || ((pixel_index2 >= 3969) && (pixel_index2 <= 3972)) || ((pixel_index2 >= 3974) && (pixel_index2 <= 3977)) || pixel_index2 == 3979 || ((pixel_index2 >= 3981) && (pixel_index2 <= 3982)) || ((pixel_index2 >= 3984) && (pixel_index2 <= 3986)) || ((pixel_index2 >= 4034) && (pixel_index2 <= 4035)) || ((pixel_index2 >= 4039) && (pixel_index2 <= 4040)) || ((pixel_index2 >= 4045) && (pixel_index2 <= 4046)) || pixel_index2 == 4048 || ((pixel_index2 >= 4050) && (pixel_index2 <= 4051)) || ((pixel_index2 >= 4057) && (pixel_index2 <= 4058)) || ((pixel_index2 >= 4060) && (pixel_index2 <= 4061)) || pixel_index2 == 4065 || ((pixel_index2 >= 4067) && (pixel_index2 <= 4068)) || pixel_index2 == 4070 || ((pixel_index2 >= 4072) && (pixel_index2 <= 4073)) || ((pixel_index2 >= 4075) && (pixel_index2 <= 4078)) || ((pixel_index2 >= 4082) && (pixel_index2 <= 4083)) || ((pixel_index2 >= 4130) && (pixel_index2 <= 4131)) || ((pixel_index2 >= 4135) && (pixel_index2 <= 4136)) || ((pixel_index2 >= 4139) && (pixel_index2 <= 4140)) || pixel_index2 == 4142 || pixel_index2 == 4144 || ((pixel_index2 >= 4146) && (pixel_index2 <= 4147)) || ((pixel_index2 >= 4151) && (pixel_index2 <= 4152)) || pixel_index2 == 4154 || ((pixel_index2 >= 4157) && (pixel_index2 <= 4159)) || pixel_index2 == 4161 || ((pixel_index2 >= 4163) && (pixel_index2 <= 4164)) || pixel_index2 == 4166 || ((pixel_index2 >= 4168) && (pixel_index2 <= 4169)) || pixel_index2 == 4171 || ((pixel_index2 >= 4173) && (pixel_index2 <= 4174)) || ((pixel_index2 >= 4178) && (pixel_index2 <= 4179)) || ((pixel_index2 >= 4225) && (pixel_index2 <= 4228)) || pixel_index2 == 4230 || pixel_index2 == 4233 || ((pixel_index2 >= 4235) && (pixel_index2 <= 4238)) || ((pixel_index2 >= 4240) && (pixel_index2 <= 4243)) || ((pixel_index2 >= 4247) && (pixel_index2 <= 4250)) || ((pixel_index2 >= 4252) && (pixel_index2 <= 4254)) || ((pixel_index2 >= 4257) && (pixel_index2 <= 4260)) || ((pixel_index2 >= 4262) && (pixel_index2 <= 4265)) || pixel_index2 == 4267 || ((pixel_index2 >= 4269) && (pixel_index2 <= 4270)) || ((pixel_index2 >= 4272) && (pixel_index2 <= 4274)) || pixel_index2 == 4802 || pixel_index2 == 4893 || pixel_index2 == 5762 || pixel_index2 == 5853) oled_data2 = 16'b1111011110011110;
                    else if (pixel_index2 == 124 || ((pixel_index2 >= 130) && (pixel_index2 <= 184)) || pixel_index2 == 190 || pixel_index2 == 220 || pixel_index2 == 229 || pixel_index2 == 233 || pixel_index2 == 237 || pixel_index2 == 241 || pixel_index2 == 245 || pixel_index2 == 249 || pixel_index2 == 253 || pixel_index2 == 257 || pixel_index2 == 261 || pixel_index2 == 265 || pixel_index2 == 269 || pixel_index2 == 273 || pixel_index2 == 277 || pixel_index2 == 286 || pixel_index2 == 316 || pixel_index2 == 325 || pixel_index2 == 329 || pixel_index2 == 333 || pixel_index2 == 337 || pixel_index2 == 341 || pixel_index2 == 345 || pixel_index2 == 349 || pixel_index2 == 353 || pixel_index2 == 357 || pixel_index2 == 361 || pixel_index2 == 365 || pixel_index2 == 369 || pixel_index2 == 373 || pixel_index2 == 382 || pixel_index2 == 412 || pixel_index2 == 421 || pixel_index2 == 425 || pixel_index2 == 429 || pixel_index2 == 433 || pixel_index2 == 437 || pixel_index2 == 441 || pixel_index2 == 445 || pixel_index2 == 449 || pixel_index2 == 453 || pixel_index2 == 457 || pixel_index2 == 461 || pixel_index2 == 465 || pixel_index2 == 469 || pixel_index2 == 478 || pixel_index2 == 508 || pixel_index2 == 517 || pixel_index2 == 521 || pixel_index2 == 525 || pixel_index2 == 529 || pixel_index2 == 533 || pixel_index2 == 537 || pixel_index2 == 541 || pixel_index2 == 545 || pixel_index2 == 549 || pixel_index2 == 553 || pixel_index2 == 557 || pixel_index2 == 561 || pixel_index2 == 565 || pixel_index2 == 574 || pixel_index2 == 604 || pixel_index2 == 613 || pixel_index2 == 617 || pixel_index2 == 621 || pixel_index2 == 625 || pixel_index2 == 629 || pixel_index2 == 633 || pixel_index2 == 637 || pixel_index2 == 641 || pixel_index2 == 645 || pixel_index2 == 649 || pixel_index2 == 653 || pixel_index2 == 657 || pixel_index2 == 661 || pixel_index2 == 670 || pixel_index2 == 700 || pixel_index2 == 709 || pixel_index2 == 713 || pixel_index2 == 717 || pixel_index2 == 721 || pixel_index2 == 725 || pixel_index2 == 729 || pixel_index2 == 733 || pixel_index2 == 737 || pixel_index2 == 741 || pixel_index2 == 745 || pixel_index2 == 749 || pixel_index2 == 753 || pixel_index2 == 757 || pixel_index2 == 766 || pixel_index2 == 796 || ((pixel_index2 >= 802) && (pixel_index2 <= 856)) || pixel_index2 == 862 || ((pixel_index2 >= 892) && (pixel_index2 <= 894)) || ((pixel_index2 >= 897) && (pixel_index2 <= 898)) || ((pixel_index2 >= 901) && (pixel_index2 <= 902)) || ((pixel_index2 >= 905) && (pixel_index2 <= 906)) || ((pixel_index2 >= 909) && (pixel_index2 <= 910)) || ((pixel_index2 >= 913) && (pixel_index2 <= 914)) || ((pixel_index2 >= 917) && (pixel_index2 <= 918)) || ((pixel_index2 >= 921) && (pixel_index2 <= 922)) || ((pixel_index2 >= 925) && (pixel_index2 <= 926)) || ((pixel_index2 >= 929) && (pixel_index2 <= 930)) || ((pixel_index2 >= 933) && (pixel_index2 <= 934)) || ((pixel_index2 >= 937) && (pixel_index2 <= 938)) || ((pixel_index2 >= 941) && (pixel_index2 <= 942)) || ((pixel_index2 >= 945) && (pixel_index2 <= 946)) || ((pixel_index2 >= 949) && (pixel_index2 <= 950)) || ((pixel_index2 >= 953) && (pixel_index2 <= 954)) || ((pixel_index2 >= 957) && (pixel_index2 <= 958)) || ((pixel_index2 >= 988) && (pixel_index2 <= 1054)) || ((pixel_index2 >= 1084) && (pixel_index2 <= 1085)) || ((pixel_index2 >= 1087) && (pixel_index2 <= 1089)) || ((pixel_index2 >= 1091) && (pixel_index2 <= 1093)) || ((pixel_index2 >= 1095) && (pixel_index2 <= 1097)) || ((pixel_index2 >= 1099) && (pixel_index2 <= 1101)) || ((pixel_index2 >= 1103) && (pixel_index2 <= 1105)) || ((pixel_index2 >= 1107) && (pixel_index2 <= 1109)) || ((pixel_index2 >= 1111) && (pixel_index2 <= 1113)) || ((pixel_index2 >= 1115) && (pixel_index2 <= 1117)) || ((pixel_index2 >= 1119) && (pixel_index2 <= 1121)) || ((pixel_index2 >= 1123) && (pixel_index2 <= 1125)) || ((pixel_index2 >= 1127) && (pixel_index2 <= 1129)) || ((pixel_index2 >= 1131) && (pixel_index2 <= 1133)) || ((pixel_index2 >= 1135) && (pixel_index2 <= 1137)) || ((pixel_index2 >= 1139) && (pixel_index2 <= 1141)) || ((pixel_index2 >= 1143) && (pixel_index2 <= 1145)) || ((pixel_index2 >= 1147) && (pixel_index2 <= 1150)) || ((pixel_index2 >= 1182) && (pixel_index2 <= 1219)) || ((pixel_index2 >= 1240) && (pixel_index2 <= 1244)) || ((pixel_index2 >= 1278) && (pixel_index2 <= 1280)) || ((pixel_index2 >= 1283) && (pixel_index2 <= 1286)) || ((pixel_index2 >= 1290) && (pixel_index2 <= 1291)) || ((pixel_index2 >= 1293) && (pixel_index2 <= 1294)) || ((pixel_index2 >= 1314) && (pixel_index2 <= 1315)) || ((pixel_index2 >= 1336) && (pixel_index2 <= 1340)) || ((pixel_index2 >= 1374) && (pixel_index2 <= 1376)) || ((pixel_index2 >= 1378) && (pixel_index2 <= 1382)) || ((pixel_index2 >= 1386) && (pixel_index2 <= 1390)) || ((pixel_index2 >= 1410) && (pixel_index2 <= 1411)) || ((pixel_index2 >= 1432) && (pixel_index2 <= 1436)) || ((pixel_index2 >= 1470) && (pixel_index2 <= 1478)) || ((pixel_index2 >= 1482) && (pixel_index2 <= 1486)) || ((pixel_index2 >= 1506) && (pixel_index2 <= 1507)) || ((pixel_index2 >= 1528) && (pixel_index2 <= 1532)) || ((pixel_index2 >= 1566) && (pixel_index2 <= 1603)) || ((pixel_index2 >= 1624) && (pixel_index2 <= 1628)) || ((pixel_index2 >= 1662) && (pixel_index2 <= 1666)) || pixel_index2 == 1670 || pixel_index2 == 1674 || ((pixel_index2 >= 1678) && (pixel_index2 <= 1696)) || ((pixel_index2 >= 1698) && (pixel_index2 <= 1699)) || ((pixel_index2 >= 1720) && (pixel_index2 <= 1724)) || ((pixel_index2 >= 1758) && (pixel_index2 <= 1762)) || pixel_index2 == 1766 || pixel_index2 == 1770 || ((pixel_index2 >= 1774) && (pixel_index2 <= 1775)) || ((pixel_index2 >= 1777) && (pixel_index2 <= 1789)) || pixel_index2 == 1792 || ((pixel_index2 >= 1794) && (pixel_index2 <= 1795)) || pixel_index2 == 1816 || ((pixel_index2 >= 1818) && (pixel_index2 <= 1820)) || ((pixel_index2 >= 1854) && (pixel_index2 <= 1858)) || pixel_index2 == 1862 || pixel_index2 == 1866 || pixel_index2 == 1870 || ((pixel_index2 >= 1872) && (pixel_index2 <= 1878)) || ((pixel_index2 >= 1882) && (pixel_index2 <= 1888)) || ((pixel_index2 >= 1892) && (pixel_index2 <= 1913)) || ((pixel_index2 >= 1915) && (pixel_index2 <= 1916)) || ((pixel_index2 >= 1948) && (pixel_index2 <= 1957)) || ((pixel_index2 >= 1963) && (pixel_index2 <= 1973)) || pixel_index2 == 1988 || pixel_index2 == 1991 || ((pixel_index2 >= 1993) && (pixel_index2 <= 1994)) || pixel_index2 == 1996 || ((pixel_index2 >= 2000) && (pixel_index2 <= 2001)) || pixel_index2 == 2008 || ((pixel_index2 >= 2011) && (pixel_index2 <= 2014)) || ((pixel_index2 >= 2044) && (pixel_index2 <= 2046)) || ((pixel_index2 >= 2048) && (pixel_index2 <= 2053)) || ((pixel_index2 >= 2059) && (pixel_index2 <= 2069)) || ((pixel_index2 >= 2084) && (pixel_index2 <= 2085)) || pixel_index2 == 2089 || ((pixel_index2 >= 2091) && (pixel_index2 <= 2093)) || ((pixel_index2 >= 2095) && (pixel_index2 <= 2096)) || ((pixel_index2 >= 2104) && (pixel_index2 <= 2105)) || ((pixel_index2 >= 2107) && (pixel_index2 <= 2110)) || pixel_index2 == 2140 || pixel_index2 == 2142 || ((pixel_index2 >= 2144) && (pixel_index2 <= 2149)) || ((pixel_index2 >= 2157) && (pixel_index2 <= 2168)) || pixel_index2 == 2178 || ((pixel_index2 >= 2180) && (pixel_index2 <= 2184)) || pixel_index2 == 2188 || ((pixel_index2 >= 2190) && (pixel_index2 <= 2192)) || ((pixel_index2 >= 2195) && (pixel_index2 <= 2197)) || ((pixel_index2 >= 2200) && (pixel_index2 <= 2206)) || ((pixel_index2 >= 2236) && (pixel_index2 <= 2238)) || pixel_index2 == 2245 || ((pixel_index2 >= 2252) && (pixel_index2 <= 2264)) || ((pixel_index2 >= 2274) && (pixel_index2 <= 2288)) || ((pixel_index2 >= 2291) && (pixel_index2 <= 2293)) || ((pixel_index2 >= 2296) && (pixel_index2 <= 2302)) || ((pixel_index2 >= 2332) && (pixel_index2 <= 2334)) || pixel_index2 == 2341 || ((pixel_index2 >= 2347) && (pixel_index2 <= 2355)) || ((pixel_index2 >= 2374) && (pixel_index2 <= 2384)) || ((pixel_index2 >= 2392) && (pixel_index2 <= 2398)) || ((pixel_index2 >= 2428) && (pixel_index2 <= 2437)) || ((pixel_index2 >= 2443) && (pixel_index2 <= 2451)) || ((pixel_index2 >= 2470) && (pixel_index2 <= 2480)) || ((pixel_index2 >= 2487) && (pixel_index2 <= 2494)) || ((pixel_index2 >= 2526) && (pixel_index2 <= 2532)) || ((pixel_index2 >= 2540) && (pixel_index2 <= 2547)) || pixel_index2 == 2566 || ((pixel_index2 >= 2580) && (pixel_index2 <= 2588)) || ((pixel_index2 >= 2622) && (pixel_index2 <= 2626)) || pixel_index2 == 2636 || ((pixel_index2 >= 2639) && (pixel_index2 <= 2644)) || ((pixel_index2 >= 2647) && (pixel_index2 <= 2648)) || pixel_index2 == 2659 || ((pixel_index2 >= 2661) && (pixel_index2 <= 2662)) || ((pixel_index2 >= 2676) && (pixel_index2 <= 2684)) || ((pixel_index2 >= 2718) && (pixel_index2 <= 2721)) || pixel_index2 == 2732 || ((pixel_index2 >= 2735) && (pixel_index2 <= 2742)) || ((pixel_index2 >= 2756) && (pixel_index2 <= 2758)) || ((pixel_index2 >= 2772) && (pixel_index2 <= 2780)) || ((pixel_index2 >= 2814) && (pixel_index2 <= 2817)) || pixel_index2 == 2828 || ((pixel_index2 >= 2831) && (pixel_index2 <= 2838)) || ((pixel_index2 >= 2842) && (pixel_index2 <= 2848)) || ((pixel_index2 >= 2852) && (pixel_index2 <= 2859)) || ((pixel_index2 >= 2866) && (pixel_index2 <= 2876)) || ((pixel_index2 >= 2910) && (pixel_index2 <= 2913)) || pixel_index2 == 2924 || ((pixel_index2 >= 2927) && (pixel_index2 <= 2935)) || ((pixel_index2 >= 2938) && (pixel_index2 <= 2944)) || ((pixel_index2 >= 2947) && (pixel_index2 <= 2955)) || pixel_index2 == 2962 || ((pixel_index2 >= 2964) && (pixel_index2 <= 2972)) || ((pixel_index2 >= 3006) && (pixel_index2 <= 3013)) || ((pixel_index2 >= 3019) && (pixel_index2 <= 3021)) || ((pixel_index2 >= 3023) && (pixel_index2 <= 3032)) || ((pixel_index2 >= 3042) && (pixel_index2 <= 3051)) || ((pixel_index2 >= 3058) && (pixel_index2 <= 3060)) || pixel_index2 == 3063 || ((pixel_index2 >= 3065) && (pixel_index2 <= 3068)) || ((pixel_index2 >= 3102) && (pixel_index2 <= 3104)) || pixel_index2 == 3107 || ((pixel_index2 >= 3117) && (pixel_index2 <= 3123)) || ((pixel_index2 >= 3143) && (pixel_index2 <= 3147)) || ((pixel_index2 >= 3154) && (pixel_index2 <= 3155)) || pixel_index2 == 3159 || ((pixel_index2 >= 3161) && (pixel_index2 <= 3164)) || ((pixel_index2 >= 3198) && (pixel_index2 <= 3200)) || ((pixel_index2 >= 3202) && (pixel_index2 <= 3203)) || ((pixel_index2 >= 3213) && (pixel_index2 <= 3216)) || ((pixel_index2 >= 3218) && (pixel_index2 <= 3219)) || ((pixel_index2 >= 3239) && (pixel_index2 <= 3243)) || ((pixel_index2 >= 3250) && (pixel_index2 <= 3251)) || ((pixel_index2 >= 3255) && (pixel_index2 <= 3260)) || ((pixel_index2 >= 3292) && (pixel_index2 <= 3299)) || ((pixel_index2 >= 3309) && (pixel_index2 <= 3312)) || ((pixel_index2 >= 3314) && (pixel_index2 <= 3315)) || ((pixel_index2 >= 3335) && (pixel_index2 <= 3337)) || pixel_index2 == 3339 || ((pixel_index2 >= 3346) && (pixel_index2 <= 3347)) || ((pixel_index2 >= 3351) && (pixel_index2 <= 3352)) || ((pixel_index2 >= 3354) && (pixel_index2 <= 3358)) || ((pixel_index2 >= 3388) && (pixel_index2 <= 3393)) || pixel_index2 == 3395 || ((pixel_index2 >= 3405) && (pixel_index2 <= 3407)) || ((pixel_index2 >= 3409) && (pixel_index2 <= 3411)) || ((pixel_index2 >= 3431) && (pixel_index2 <= 3432)) || ((pixel_index2 >= 3434) && (pixel_index2 <= 3435)) || ((pixel_index2 >= 3438) && (pixel_index2 <= 3443)) || ((pixel_index2 >= 3447) && (pixel_index2 <= 3448)) || ((pixel_index2 >= 3450) && (pixel_index2 <= 3454)) || ((pixel_index2 >= 3484) && (pixel_index2 <= 3487)) || pixel_index2 == 3489 || pixel_index2 == 3491 || ((pixel_index2 >= 3501) && (pixel_index2 <= 3502)) || ((pixel_index2 >= 3505) && (pixel_index2 <= 3507)) || ((pixel_index2 >= 3527) && (pixel_index2 <= 3531)) || ((pixel_index2 >= 3538) && (pixel_index2 <= 3539)) || ((pixel_index2 >= 3543) && (pixel_index2 <= 3544)) || ((pixel_index2 >= 3546) && (pixel_index2 <= 3550)) || ((pixel_index2 >= 3580) && (pixel_index2 <= 3587)) || ((pixel_index2 >= 3597) && (pixel_index2 <= 3603)) || ((pixel_index2 >= 3623) && (pixel_index2 <= 3628)) || ((pixel_index2 >= 3633) && (pixel_index2 <= 3635)) || ((pixel_index2 >= 3639) && (pixel_index2 <= 3646)) || ((pixel_index2 >= 4620) && (pixel_index2 <= 4692)) || ((pixel_index2 >= 4707) && (pixel_index2 <= 4796)) || ((pixel_index2 >= 4803) && (pixel_index2 <= 4812)) || ((pixel_index2 >= 4814) && (pixel_index2 <= 4817)) || ((pixel_index2 >= 4819) && (pixel_index2 <= 4820)) || ((pixel_index2 >= 4827) && (pixel_index2 <= 4829)) || ((pixel_index2 >= 4834) && (pixel_index2 <= 4835)) || ((pixel_index2 >= 4838) && (pixel_index2 <= 4839)) || ((pixel_index2 >= 4841) && (pixel_index2 <= 4843)) || ((pixel_index2 >= 4845) && (pixel_index2 <= 4846)) || ((pixel_index2 >= 4851) && (pixel_index2 <= 4861)) || ((pixel_index2 >= 4863) && (pixel_index2 <= 4865)) || ((pixel_index2 >= 4868) && (pixel_index2 <= 4869)) || ((pixel_index2 >= 4871) && (pixel_index2 <= 4873)) || ((pixel_index2 >= 4880) && (pixel_index2 <= 4882)) || ((pixel_index2 >= 4887) && (pixel_index2 <= 4892)) || ((pixel_index2 >= 4899) && (pixel_index2 <= 4907)) || ((pixel_index2 >= 4910) && (pixel_index2 <= 4912)) || pixel_index2 == 4915 || pixel_index2 == 4924 || pixel_index2 == 4931 || pixel_index2 == 4935 || pixel_index2 == 4938 || pixel_index2 == 4941 || ((pixel_index2 >= 4948) && (pixel_index2 <= 4956)) || ((pixel_index2 >= 4959) && (pixel_index2 <= 4961)) || pixel_index2 == 4965 || pixel_index2 == 4968 || pixel_index2 == 4977 || ((pixel_index2 >= 4984) && (pixel_index2 <= 4988)) || ((pixel_index2 >= 4994) && (pixel_index2 <= 5003)) || ((pixel_index2 >= 5006) && (pixel_index2 <= 5008)) || pixel_index2 == 5011 || pixel_index2 == 5020 || pixel_index2 == 5027 || pixel_index2 == 5034 || pixel_index2 == 5037 || ((pixel_index2 >= 5044) && (pixel_index2 <= 5052)) || ((pixel_index2 >= 5055) && (pixel_index2 <= 5057)) || pixel_index2 == 5064 || pixel_index2 == 5073 || ((pixel_index2 >= 5080) && (pixel_index2 <= 5085)) || ((pixel_index2 >= 5090) && (pixel_index2 <= 5099)) || ((pixel_index2 >= 5102) && (pixel_index2 <= 5104)) || pixel_index2 == 5107 || ((pixel_index2 >= 5111) && (pixel_index2 <= 5112)) || ((pixel_index2 >= 5116) && (pixel_index2 <= 5119)) || ((pixel_index2 >= 5123) && (pixel_index2 <= 5124)) || pixel_index2 == 5130 || ((pixel_index2 >= 5133) && (pixel_index2 <= 5136)) || ((pixel_index2 >= 5140) && (pixel_index2 <= 5148)) || ((pixel_index2 >= 5151) && (pixel_index2 <= 5154)) || pixel_index2 == 5160 || ((pixel_index2 >= 5164) && (pixel_index2 <= 5165)) || pixel_index2 == 5169 || ((pixel_index2 >= 5173) && (pixel_index2 <= 5181)) || ((pixel_index2 >= 5186) && (pixel_index2 <= 5195)) || ((pixel_index2 >= 5198) && (pixel_index2 <= 5200)) || pixel_index2 == 5203 || ((pixel_index2 >= 5206) && (pixel_index2 <= 5209)) || ((pixel_index2 >= 5212) && (pixel_index2 <= 5216)) || ((pixel_index2 >= 5219) && (pixel_index2 <= 5220)) || pixel_index2 == 5226 || ((pixel_index2 >= 5229) && (pixel_index2 <= 5233)) || ((pixel_index2 >= 5236) && (pixel_index2 <= 5244)) || ((pixel_index2 >= 5247) && (pixel_index2 <= 5250)) || pixel_index2 == 5256 || ((pixel_index2 >= 5259) && (pixel_index2 <= 5262)) || pixel_index2 == 5265 || ((pixel_index2 >= 5271) && (pixel_index2 <= 5277)) || ((pixel_index2 >= 5282) && (pixel_index2 <= 5291)) || ((pixel_index2 >= 5294) && (pixel_index2 <= 5296)) || pixel_index2 == 5299 || ((pixel_index2 >= 5302) && (pixel_index2 <= 5305)) || ((pixel_index2 >= 5308) && (pixel_index2 <= 5312)) || pixel_index2 == 5315 || pixel_index2 == 5322 || ((pixel_index2 >= 5325) && (pixel_index2 <= 5329)) || ((pixel_index2 >= 5332) && (pixel_index2 <= 5340)) || ((pixel_index2 >= 5343) && (pixel_index2 <= 5345)) || pixel_index2 == 5352 || ((pixel_index2 >= 5355) && (pixel_index2 <= 5358)) || pixel_index2 == 5361 || ((pixel_index2 >= 5368) && (pixel_index2 <= 5373)) || ((pixel_index2 >= 5378) && (pixel_index2 <= 5387)) || ((pixel_index2 >= 5390) && (pixel_index2 <= 5392)) || pixel_index2 == 5395 || ((pixel_index2 >= 5398) && (pixel_index2 <= 5401)) || ((pixel_index2 >= 5404) && (pixel_index2 <= 5408)) || pixel_index2 == 5411 || pixel_index2 == 5415 || pixel_index2 == 5418 || ((pixel_index2 >= 5421) && (pixel_index2 <= 5425)) || ((pixel_index2 >= 5428) && (pixel_index2 <= 5436)) || ((pixel_index2 >= 5439) && (pixel_index2 <= 5441)) || pixel_index2 == 5445 || pixel_index2 == 5448 || ((pixel_index2 >= 5451) && (pixel_index2 <= 5454)) || ((pixel_index2 >= 5457) && (pixel_index2 <= 5458)) || ((pixel_index2 >= 5464) && (pixel_index2 <= 5469)) || ((pixel_index2 >= 5474) && (pixel_index2 <= 5483)) || ((pixel_index2 >= 5486) && (pixel_index2 <= 5488)) || pixel_index2 == 5491 || ((pixel_index2 >= 5494) && (pixel_index2 <= 5497)) || ((pixel_index2 >= 5500) && (pixel_index2 <= 5503)) || pixel_index2 == 5507 || ((pixel_index2 >= 5510) && (pixel_index2 <= 5511)) || pixel_index2 == 5514 || ((pixel_index2 >= 5517) && (pixel_index2 <= 5520)) || ((pixel_index2 >= 5524) && (pixel_index2 <= 5532)) || ((pixel_index2 >= 5535) && (pixel_index2 <= 5537)) || ((pixel_index2 >= 5540) && (pixel_index2 <= 5541)) || pixel_index2 == 5544 || ((pixel_index2 >= 5548) && (pixel_index2 <= 5549)) || ((pixel_index2 >= 5553) && (pixel_index2 <= 5556)) || ((pixel_index2 >= 5560) && (pixel_index2 <= 5565)) || ((pixel_index2 >= 5570) && (pixel_index2 <= 5575)) || pixel_index2 == 5584 || pixel_index2 == 5587 || ((pixel_index2 >= 5590) && (pixel_index2 <= 5593)) || pixel_index2 == 5596 || pixel_index2 == 5603 || pixel_index2 == 5610 || pixel_index2 == 5613 || ((pixel_index2 >= 5620) && (pixel_index2 <= 5624)) || pixel_index2 == 5633 || pixel_index2 == 5640 || pixel_index2 == 5649 || ((pixel_index2 >= 5656) && (pixel_index2 <= 5661)) || ((pixel_index2 >= 5667) && (pixel_index2 <= 5671)) || pixel_index2 == 5680 || pixel_index2 == 5683 || ((pixel_index2 >= 5686) && (pixel_index2 <= 5689)) || pixel_index2 == 5692 || pixel_index2 == 5699 || pixel_index2 == 5706 || pixel_index2 == 5709 || ((pixel_index2 >= 5716) && (pixel_index2 <= 5720)) || pixel_index2 == 5729 || pixel_index2 == 5736 || pixel_index2 == 5745 || ((pixel_index2 >= 5752) && (pixel_index2 <= 5756)) || ((pixel_index2 >= 5763) && (pixel_index2 <= 5768)) || ((pixel_index2 >= 5775) && (pixel_index2 <= 5776)) || ((pixel_index2 >= 5778) && (pixel_index2 <= 5780)) || ((pixel_index2 >= 5782) && (pixel_index2 <= 5785)) || ((pixel_index2 >= 5787) && (pixel_index2 <= 5789)) || ((pixel_index2 >= 5794) && (pixel_index2 <= 5796)) || ((pixel_index2 >= 5801) && (pixel_index2 <= 5802)) || ((pixel_index2 >= 5804) && (pixel_index2 <= 5806)) || ((pixel_index2 >= 5811) && (pixel_index2 <= 5817)) || ((pixel_index2 >= 5824) && (pixel_index2 <= 5826)) || ((pixel_index2 >= 5831) && (pixel_index2 <= 5833)) || ((pixel_index2 >= 5840) && (pixel_index2 <= 5842)) || ((pixel_index2 >= 5847) && (pixel_index2 <= 5852)) || (pixel_index2 >= 5868) && (pixel_index2 <= 5940)) oled_data2 = 16'b0000000000001010;
                    else if (((pixel_index2 >= 125) && (pixel_index2 <= 129)) || pixel_index2 == 221 || pixel_index2 == 225 || pixel_index2 == 317 || pixel_index2 == 321 || pixel_index2 == 413 || pixel_index2 == 417 || pixel_index2 == 509 || pixel_index2 == 513 || pixel_index2 == 605 || pixel_index2 == 609 || pixel_index2 == 701 || pixel_index2 == 705 || ((pixel_index2 >= 797) && (pixel_index2 <= 801)) || pixel_index2 == 1155 || ((pixel_index2 >= 1159) && (pixel_index2 <= 1161)) || pixel_index2 == 1163 || ((pixel_index2 >= 1165) && (pixel_index2 <= 1166)) || pixel_index2 == 1168 || ((pixel_index2 >= 1170) && (pixel_index2 <= 1171)) || pixel_index2 == 1173 || ((pixel_index2 >= 1175) && (pixel_index2 <= 1176)) || pixel_index2 == 1178 || pixel_index2 == 1254 || ((pixel_index2 >= 1256) && (pixel_index2 <= 1257)) || pixel_index2 == 1259 || ((pixel_index2 >= 1261) && (pixel_index2 <= 1262)) || ((pixel_index2 >= 1264) && (pixel_index2 <= 1267)) || ((pixel_index2 >= 1270) && (pixel_index2 <= 1272)) || pixel_index2 == 1350 || ((pixel_index2 >= 1352) && (pixel_index2 <= 1353)) || pixel_index2 == 1355 || ((pixel_index2 >= 1357) && (pixel_index2 <= 1358)) || pixel_index2 == 1360 || ((pixel_index2 >= 1362) && (pixel_index2 <= 1363)) || pixel_index2 == 1365 || ((pixel_index2 >= 1367) && (pixel_index2 <= 1368)) || ((pixel_index2 >= 1447) && (pixel_index2 <= 1449)) || ((pixel_index2 >= 1451) && (pixel_index2 <= 1454)) || ((pixel_index2 >= 1456) && (pixel_index2 <= 1459)) || ((pixel_index2 >= 1461) && (pixel_index2 <= 1464)) || pixel_index2 == 1466) oled_data2 = 16'b1010001010010100;
                    else if (((pixel_index2 >= 185) && (pixel_index2 <= 189)) || pixel_index2 == 281 || pixel_index2 == 285 || pixel_index2 == 377 || pixel_index2 == 381 || pixel_index2 == 473 || pixel_index2 == 477 || pixel_index2 == 569 || pixel_index2 == 573 || pixel_index2 == 665 || pixel_index2 == 669 || pixel_index2 == 761 || pixel_index2 == 765 || ((pixel_index2 >= 857) && (pixel_index2 <= 861)) || ((pixel_index2 >= 4008) && (pixel_index2 <= 4009)) || ((pixel_index2 >= 4012) && (pixel_index2 <= 4015)) || ((pixel_index2 >= 4017) && (pixel_index2 <= 4020)) || ((pixel_index2 >= 4022) && (pixel_index2 <= 4025)) || pixel_index2 == 4027 || ((pixel_index2 >= 4029) && (pixel_index2 <= 4030)) || ((pixel_index2 >= 4104) && (pixel_index2 <= 4105)) || ((pixel_index2 >= 4110) && (pixel_index2 <= 4111)) || ((pixel_index2 >= 4113) && (pixel_index2 <= 4114)) || ((pixel_index2 >= 4120) && (pixel_index2 <= 4121)) || ((pixel_index2 >= 4124) && (pixel_index2 <= 4126)) || ((pixel_index2 >= 4200) && (pixel_index2 <= 4201)) || ((pixel_index2 >= 4204) && (pixel_index2 <= 4205)) || pixel_index2 == 4207 || ((pixel_index2 >= 4210) && (pixel_index2 <= 4212)) || ((pixel_index2 >= 4214) && (pixel_index2 <= 4215)) || pixel_index2 == 4217 || pixel_index2 == 4219 || ((pixel_index2 >= 4221) && (pixel_index2 <= 4222)) || ((pixel_index2 >= 4295) && (pixel_index2 <= 4298)) || ((pixel_index2 >= 4300) && (pixel_index2 <= 4303)) || ((pixel_index2 >= 4305) && (pixel_index2 <= 4307)) || ((pixel_index2 >= 4310) && (pixel_index2 <= 4313)) || (pixel_index2 >= 4315) && (pixel_index2 <= 4318)) oled_data2 = 16'b0101011110010100;
                    else if (pixel_index2 == 319 || pixel_index2 == 331 || pixel_index2 == 335 || pixel_index2 == 339 || pixel_index2 == 343 || pixel_index2 == 347 || pixel_index2 == 415 || pixel_index2 == 427 || pixel_index2 == 431 || pixel_index2 == 435 || pixel_index2 == 439 || pixel_index2 == 443 || pixel_index2 == 3253 || pixel_index2 == 3349) oled_data2 = 16'b0000010100000000;
                    else if (pixel_index2 == 515 || pixel_index2 == 519 || pixel_index2 == 543 || pixel_index2 == 547 || pixel_index2 == 551 || pixel_index2 == 555 || pixel_index2 == 559 || pixel_index2 == 563 || pixel_index2 == 567 || pixel_index2 == 571 || pixel_index2 == 611 || pixel_index2 == 615 || pixel_index2 == 639 || pixel_index2 == 643 || pixel_index2 == 647 || pixel_index2 == 651 || pixel_index2 == 655 || pixel_index2 == 659 || pixel_index2 == 663 || pixel_index2 == 667 || pixel_index2 == 3488) oled_data2 = 16'b1010000000000000;
                    else if (pixel_index2 == 1086 || pixel_index2 == 1090 || pixel_index2 == 1094 || pixel_index2 == 1118 || pixel_index2 == 1122 || pixel_index2 == 1126 || pixel_index2 == 1130 || pixel_index2 == 1134 || pixel_index2 == 1138 || pixel_index2 == 1142 || pixel_index2 == 1146) oled_data2 = 16'b0000001010000000;
                    else if (pixel_index2 == 1098 || pixel_index2 == 1102 || pixel_index2 == 1106 || pixel_index2 == 1110 || pixel_index2 == 1114) oled_data2 = 16'b1111011110001010;
                    else if (((pixel_index2 >= 1281) && (pixel_index2 <= 1282)) || pixel_index2 == 1292 || pixel_index2 == 1295 || ((pixel_index2 >= 1297) && (pixel_index2 <= 1299)) || pixel_index2 == 1302 || ((pixel_index2 >= 1304) && (pixel_index2 <= 1305)) || pixel_index2 == 1307 || pixel_index2 == 1309 || pixel_index2 == 1311 || pixel_index2 == 1313 || pixel_index2 == 1377 || ((pixel_index2 >= 1392) && (pixel_index2 <= 1395)) || ((pixel_index2 >= 1397) && (pixel_index2 <= 1399)) || pixel_index2 == 1401 || ((pixel_index2 >= 1403) && (pixel_index2 <= 1404)) || pixel_index2 == 1406 || pixel_index2 == 1409 || ((pixel_index2 >= 1487) && (pixel_index2 <= 1488)) || pixel_index2 == 1490 || pixel_index2 == 1493 || pixel_index2 == 1495 || pixel_index2 == 1497 || ((pixel_index2 >= 1499) && (pixel_index2 <= 1500)) || ((pixel_index2 >= 1502) && (pixel_index2 <= 1503)) || pixel_index2 == 1505 || pixel_index2 == 1697 || pixel_index2 == 1776 || ((pixel_index2 >= 1790) && (pixel_index2 <= 1791)) || pixel_index2 == 1793 || pixel_index2 == 1817 || pixel_index2 == 1871 || pixel_index2 == 1914 || pixel_index2 == 1974 || ((pixel_index2 >= 1989) && (pixel_index2 <= 1990)) || pixel_index2 == 1992 || pixel_index2 == 1995 || ((pixel_index2 >= 1997) && (pixel_index2 <= 1999)) || ((pixel_index2 >= 2009) && (pixel_index2 <= 2010)) || pixel_index2 == 2047 || ((pixel_index2 >= 2070) && (pixel_index2 <= 2071)) || pixel_index2 == 2083 || ((pixel_index2 >= 2086) && (pixel_index2 <= 2088)) || pixel_index2 == 2090 || pixel_index2 == 2094 || pixel_index2 == 2106 || pixel_index2 == 2141 || pixel_index2 == 2143 || ((pixel_index2 >= 2155) && (pixel_index2 <= 2156)) || pixel_index2 == 2179 || ((pixel_index2 >= 2185) && (pixel_index2 <= 2187)) || pixel_index2 == 2189 || pixel_index2 == 2240 || pixel_index2 == 2243 || pixel_index2 == 2251 || pixel_index2 == 2336 || pixel_index2 == 2338 || pixel_index2 == 2340 || pixel_index2 == 2548 || ((pixel_index2 >= 2550) && (pixel_index2 <= 2551)) || ((pixel_index2 >= 2562) && (pixel_index2 <= 2563)) || ((pixel_index2 >= 2567) && (pixel_index2 <= 2579)) || ((pixel_index2 >= 2645) && (pixel_index2 <= 2646)) || pixel_index2 == 2658 || pixel_index2 == 2660 || ((pixel_index2 >= 2663) && (pixel_index2 <= 2675)) || ((pixel_index2 >= 2759) && (pixel_index2 <= 2771)) || ((pixel_index2 >= 2925) && (pixel_index2 <= 2926)) || pixel_index2 == 2937 || pixel_index2 == 2946 || pixel_index2 == 3022 || ((pixel_index2 >= 3105) && (pixel_index2 <= 3106)) || pixel_index2 == 3201 || pixel_index2 == 3217 || ((pixel_index2 >= 3230) && (pixel_index2 <= 3231)) || pixel_index2 == 3313 || pixel_index2 == 3324 || pixel_index2 == 3408 || ((pixel_index2 >= 3421) && (pixel_index2 <= 3422)) || ((pixel_index2 >= 3503) && (pixel_index2 <= 3504)) || ((pixel_index2 >= 3533) && (pixel_index2 <= 3536)) || pixel_index2 == 3629 || pixel_index2 == 3632) oled_data2 = 16'b1010010100010100;
                    else if (pixel_index2 == 1287 || pixel_index2 == 1289 || pixel_index2 == 1479 || pixel_index2 == 1481 || pixel_index2 == 1667 || pixel_index2 == 1669 || pixel_index2 == 1671 || pixel_index2 == 1673 || pixel_index2 == 1675 || pixel_index2 == 1677 || pixel_index2 == 1859 || pixel_index2 == 1861 || pixel_index2 == 1863 || pixel_index2 == 1865 || pixel_index2 == 1867 || pixel_index2 == 1869 || ((pixel_index2 >= 1879) && (pixel_index2 <= 1881)) || ((pixel_index2 >= 1889) && (pixel_index2 <= 1891)) || ((pixel_index2 >= 1975) && (pixel_index2 <= 1987)) || ((pixel_index2 >= 2002) && (pixel_index2 <= 2007)) || pixel_index2 == 2055 || pixel_index2 == 2057 || ((pixel_index2 >= 2072) && (pixel_index2 <= 2073)) || ((pixel_index2 >= 2081) && (pixel_index2 <= 2082)) || ((pixel_index2 >= 2097) && (pixel_index2 <= 2103)) || pixel_index2 == 2169 || pixel_index2 == 2177 || ((pixel_index2 >= 2193) && (pixel_index2 <= 2194)) || ((pixel_index2 >= 2198) && (pixel_index2 <= 2199)) || pixel_index2 == 2239 || ((pixel_index2 >= 2241) && (pixel_index2 <= 2242)) || pixel_index2 == 2244 || pixel_index2 == 2247 || pixel_index2 == 2249 || pixel_index2 == 2265 || pixel_index2 == 2273 || ((pixel_index2 >= 2289) && (pixel_index2 <= 2290)) || ((pixel_index2 >= 2294) && (pixel_index2 <= 2295)) || pixel_index2 == 2335 || pixel_index2 == 2337 || pixel_index2 == 2339 || ((pixel_index2 >= 2356) && (pixel_index2 <= 2361)) || ((pixel_index2 >= 2369) && (pixel_index2 <= 2373)) || ((pixel_index2 >= 2385) && (pixel_index2 <= 2391)) || ((pixel_index2 >= 2438) && (pixel_index2 <= 2442)) || ((pixel_index2 >= 2452) && (pixel_index2 <= 2457)) || ((pixel_index2 >= 2465) && (pixel_index2 <= 2469)) || ((pixel_index2 >= 2481) && (pixel_index2 <= 2486)) || pixel_index2 == 2533 || pixel_index2 == 2539 || pixel_index2 == 2549 || ((pixel_index2 >= 2552) && (pixel_index2 <= 2553)) || pixel_index2 == 2561 || ((pixel_index2 >= 2564) && (pixel_index2 <= 2565)) || ((pixel_index2 >= 2627) && (pixel_index2 <= 2629)) || pixel_index2 == 2635 || ((pixel_index2 >= 2637) && (pixel_index2 <= 2638)) || pixel_index2 == 2649 || pixel_index2 == 2657 || ((pixel_index2 >= 2722) && (pixel_index2 <= 2725)) || pixel_index2 == 2731 || ((pixel_index2 >= 2733) && (pixel_index2 <= 2734)) || ((pixel_index2 >= 2743) && (pixel_index2 <= 2755)) || ((pixel_index2 >= 2818) && (pixel_index2 <= 2821)) || pixel_index2 == 2827 || ((pixel_index2 >= 2829) && (pixel_index2 <= 2830)) || ((pixel_index2 >= 2839) && (pixel_index2 <= 2841)) || ((pixel_index2 >= 2849) && (pixel_index2 <= 2851)) || ((pixel_index2 >= 2914) && (pixel_index2 <= 2917)) || pixel_index2 == 2923 || pixel_index2 == 2936 || pixel_index2 == 2945 || pixel_index2 == 2963 || ((pixel_index2 >= 3014) && (pixel_index2 <= 3018)) || ((pixel_index2 >= 3061) && (pixel_index2 <= 3062)) || pixel_index2 == 3064 || ((pixel_index2 >= 3108) && (pixel_index2 <= 3116)) || pixel_index2 == 3160 || ((pixel_index2 >= 3204) && (pixel_index2 <= 3212)) || ((pixel_index2 >= 3300) && (pixel_index2 <= 3308)) || pixel_index2 == 3317 || ((pixel_index2 >= 3319) && (pixel_index2 <= 3320)) || ((pixel_index2 >= 3330) && (pixel_index2 <= 3331)) || pixel_index2 == 3333 || pixel_index2 == 3338 || ((pixel_index2 >= 3396) && (pixel_index2 <= 3404)) || pixel_index2 == 3433 || ((pixel_index2 >= 3436) && (pixel_index2 <= 3437)) || ((pixel_index2 >= 3492) && (pixel_index2 <= 3500)) || ((pixel_index2 >= 3588) && (pixel_index2 <= 3596)) || ((pixel_index2 >= 3684) && (pixel_index2 <= 3692)) || ((pixel_index2 >= 3724) && (pixel_index2 <= 3729)) || ((pixel_index2 >= 3820) && (pixel_index2 <= 3825)) || ((pixel_index2 >= 3893) && (pixel_index2 <= 3894)) || ((pixel_index2 >= 3897) && (pixel_index2 <= 3905)) || ((pixel_index2 >= 3908) && (pixel_index2 <= 3909)) || ((pixel_index2 >= 3989) && (pixel_index2 <= 3990)) || ((pixel_index2 >= 3994) && (pixel_index2 <= 4000)) || ((pixel_index2 >= 4004) && (pixel_index2 <= 4005)) || ((pixel_index2 >= 4085) && (pixel_index2 <= 4086)) || ((pixel_index2 >= 4090) && (pixel_index2 <= 4096)) || ((pixel_index2 >= 4100) && (pixel_index2 <= 4101)) || pixel_index2 == 4706 || pixel_index2 == 4797 || pixel_index2 == 5666 || pixel_index2 == 5757) oled_data2 = 16'b0101001010001010;
                    else if (pixel_index2 == 1296 || ((pixel_index2 >= 1300) && (pixel_index2 <= 1301)) || pixel_index2 == 1303 || pixel_index2 == 1306 || pixel_index2 == 1308 || pixel_index2 == 1310 || pixel_index2 == 1312 || pixel_index2 == 1391 || pixel_index2 == 1396 || pixel_index2 == 1400 || pixel_index2 == 1402 || pixel_index2 == 1405 || ((pixel_index2 >= 1407) && (pixel_index2 <= 1408)) || pixel_index2 == 1489 || ((pixel_index2 >= 1491) && (pixel_index2 <= 1492)) || pixel_index2 == 1494 || pixel_index2 == 1496 || pixel_index2 == 1498 || pixel_index2 == 1501 || pixel_index2 == 1504 || pixel_index2 == 3353 || pixel_index2 == 3449 || pixel_index2 == 3545) oled_data2 = 16'b0101001010010100;
                    else if (((pixel_index2 >= 1317) && (pixel_index2 <= 1319)) || ((pixel_index2 >= 1322) && (pixel_index2 <= 1324)) || ((pixel_index2 >= 1327) && (pixel_index2 <= 1329)) || ((pixel_index2 >= 1332) && (pixel_index2 <= 1334)) || pixel_index2 == 1415 || pixel_index2 == 1418 || pixel_index2 == 1420 || pixel_index2 == 1423 || pixel_index2 == 1425 || pixel_index2 == 1428 || pixel_index2 == 1430 || pixel_index2 == 1511 || ((pixel_index2 >= 1514) && (pixel_index2 <= 1516)) || pixel_index2 == 1519 || pixel_index2 == 1521 || ((pixel_index2 >= 1524) && (pixel_index2 <= 1526)) || pixel_index2 == 1607 || pixel_index2 == 1612 || pixel_index2 == 1615 || pixel_index2 == 1617 || pixel_index2 == 1622 || pixel_index2 == 1703 || pixel_index2 == 1708 || pixel_index2 == 1711 || pixel_index2 == 1713 || pixel_index2 == 1718) oled_data2 = 16'b1010000000001010;
                    else if (((pixel_index2 >= 1958) && (pixel_index2 <= 1962)) || pixel_index2 == 2054 || pixel_index2 == 2058 || pixel_index2 == 2150 || pixel_index2 == 2154 || pixel_index2 == 2246 || pixel_index2 == 2250 || ((pixel_index2 >= 2342) && (pixel_index2 <= 2346)) || ((pixel_index2 >= 3364) && (pixel_index2 <= 3367)) || ((pixel_index2 >= 3370) && (pixel_index2 <= 3372)) || ((pixel_index2 >= 3375) && (pixel_index2 <= 3376)) || ((pixel_index2 >= 3380) && (pixel_index2 <= 3382)) || pixel_index2 == 3463 || pixel_index2 == 3465 || pixel_index2 == 3468 || pixel_index2 == 3470 || pixel_index2 == 3473 || pixel_index2 == 3475 || pixel_index2 == 3478 || pixel_index2 == 3481 || pixel_index2 == 3559 || ((pixel_index2 >= 3562) && (pixel_index2 <= 3564)) || pixel_index2 == 3566 || pixel_index2 == 3569 || ((pixel_index2 >= 3572) && (pixel_index2 <= 3574)) || pixel_index2 == 3576 || pixel_index2 == 3655 || pixel_index2 == 3657 || pixel_index2 == 3660 || pixel_index2 == 3662 || pixel_index2 == 3665 || pixel_index2 == 3667 || pixel_index2 == 3670 || pixel_index2 == 3673 || pixel_index2 == 3751 || ((pixel_index2 >= 3754) && (pixel_index2 <= 3756)) || pixel_index2 == 3758 || pixel_index2 == 3761 || (pixel_index2 >= 3764) && (pixel_index2 <= 3766)) oled_data2 = 16'b1010001010001010;
                    else if (pixel_index2 == 3229 || (pixel_index2 >= 3325) && (pixel_index2 <= 3326)) oled_data2 = 16'b0101010100001010;
                    else if (pixel_index2 == 3394 || pixel_index2 == 3490) oled_data2 = 16'b0000000000010100;
                    else if (pixel_index2 == 3532 || pixel_index2 == 3537) oled_data2 = 16'b0101000000000000;
                    else if (((pixel_index2 >= 4423) && (pixel_index2 <= 4505)) || ((pixel_index2 >= 4513) && (pixel_index2 <= 4518)) || (pixel_index2 >= 4602) && (pixel_index2 <= 4606)) oled_data2 = 16'b0000001010011110;
                    else if (((pixel_index2 >= 4519) && (pixel_index2 <= 4601)) || ((pixel_index2 >= 4609) && (pixel_index2 <= 4619)) || ((pixel_index2 >= 4693) && (pixel_index2 <= 4702)) || pixel_index2 == 4705 || pixel_index2 == 4798 || pixel_index2 == 4801 || pixel_index2 == 4894 || ((pixel_index2 >= 4897) && (pixel_index2 <= 4898)) || ((pixel_index2 >= 4989) && (pixel_index2 <= 4990)) || pixel_index2 == 4993 || pixel_index2 == 5086 || pixel_index2 == 5089 || pixel_index2 == 5182 || pixel_index2 == 5185 || pixel_index2 == 5278 || pixel_index2 == 5281 || pixel_index2 == 5374 || pixel_index2 == 5377 || pixel_index2 == 5470 || pixel_index2 == 5473 || pixel_index2 == 5566 || pixel_index2 == 5569 || pixel_index2 == 5662 || pixel_index2 == 5665 || pixel_index2 == 5758 || pixel_index2 == 5761 || pixel_index2 == 5854 || ((pixel_index2 >= 5857) && (pixel_index2 <= 5867)) || ((pixel_index2 >= 5941) && (pixel_index2 <= 5950)) || (pixel_index2 >= 5959) && (pixel_index2 <= 6041)) oled_data2 = 16'b0000001010010100;
                    else if (pixel_index2 == 4813 || pixel_index2 == 4818 || ((pixel_index2 >= 4821) && (pixel_index2 <= 4826)) || ((pixel_index2 >= 4830) && (pixel_index2 <= 4833)) || ((pixel_index2 >= 4836) && (pixel_index2 <= 4837)) || pixel_index2 == 4840 || pixel_index2 == 4844 || ((pixel_index2 >= 4847) && (pixel_index2 <= 4850)) || pixel_index2 == 4862 || ((pixel_index2 >= 4866) && (pixel_index2 <= 4867)) || pixel_index2 == 4870 || ((pixel_index2 >= 4874) && (pixel_index2 <= 4879)) || ((pixel_index2 >= 4883) && (pixel_index2 <= 4886)) || pixel_index2 == 4908 || pixel_index2 == 4913 || pixel_index2 == 4916 || pixel_index2 == 4923 || pixel_index2 == 4925 || pixel_index2 == 4930 || pixel_index2 == 4934 || pixel_index2 == 4937 || pixel_index2 == 4939 || pixel_index2 == 4942 || pixel_index2 == 4947 || pixel_index2 == 4957 || pixel_index2 == 4964 || pixel_index2 == 4967 || pixel_index2 == 4969 || pixel_index2 == 4976 || pixel_index2 == 4978 || pixel_index2 == 4983 || pixel_index2 == 5031 || pixel_index2 == 5061 || pixel_index2 == 5221 || pixel_index2 == 5251 || ((pixel_index2 >= 5268) && (pixel_index2 <= 5270)) || pixel_index2 == 5316 || pixel_index2 == 5346 || pixel_index2 == 5367 || pixel_index2 == 5504 || pixel_index2 == 5521 || pixel_index2 == 5547 || pixel_index2 == 5550 || pixel_index2 == 5557 || ((pixel_index2 >= 5576) && (pixel_index2 <= 5579)) || ((pixel_index2 >= 5582) && (pixel_index2 <= 5583)) || ((pixel_index2 >= 5597) && (pixel_index2 <= 5599)) || ((pixel_index2 >= 5606) && (pixel_index2 <= 5607)) || ((pixel_index2 >= 5614) && (pixel_index2 <= 5616)) || ((pixel_index2 >= 5625) && (pixel_index2 <= 5628)) || ((pixel_index2 >= 5631) && (pixel_index2 <= 5632)) || ((pixel_index2 >= 5636) && (pixel_index2 <= 5637)) || ((pixel_index2 >= 5644) && (pixel_index2 <= 5645)) || (pixel_index2 >= 5650) && (pixel_index2 <= 5652)) oled_data2 = 16'b0101001010000000;
                    else if (pixel_index2 == 4909 || pixel_index2 == 4914 || ((pixel_index2 >= 4917) && (pixel_index2 <= 4922)) || ((pixel_index2 >= 4926) && (pixel_index2 <= 4929)) || ((pixel_index2 >= 4932) && (pixel_index2 <= 4933)) || pixel_index2 == 4936 || pixel_index2 == 4940 || ((pixel_index2 >= 4943) && (pixel_index2 <= 4946)) || pixel_index2 == 4958 || ((pixel_index2 >= 4962) && (pixel_index2 <= 4963)) || pixel_index2 == 4966 || ((pixel_index2 >= 4970) && (pixel_index2 <= 4975)) || ((pixel_index2 >= 4979) && (pixel_index2 <= 4982)) || ((pixel_index2 >= 5004) && (pixel_index2 <= 5005)) || ((pixel_index2 >= 5009) && (pixel_index2 <= 5010)) || ((pixel_index2 >= 5012) && (pixel_index2 <= 5019)) || ((pixel_index2 >= 5021) && (pixel_index2 <= 5026)) || ((pixel_index2 >= 5028) && (pixel_index2 <= 5030)) || ((pixel_index2 >= 5032) && (pixel_index2 <= 5033)) || ((pixel_index2 >= 5035) && (pixel_index2 <= 5036)) || ((pixel_index2 >= 5038) && (pixel_index2 <= 5043)) || ((pixel_index2 >= 5053) && (pixel_index2 <= 5054)) || ((pixel_index2 >= 5058) && (pixel_index2 <= 5060)) || ((pixel_index2 >= 5062) && (pixel_index2 <= 5063)) || ((pixel_index2 >= 5065) && (pixel_index2 <= 5072)) || ((pixel_index2 >= 5074) && (pixel_index2 <= 5079)) || ((pixel_index2 >= 5100) && (pixel_index2 <= 5101)) || ((pixel_index2 >= 5105) && (pixel_index2 <= 5106)) || ((pixel_index2 >= 5108) && (pixel_index2 <= 5110)) || ((pixel_index2 >= 5113) && (pixel_index2 <= 5115)) || ((pixel_index2 >= 5120) && (pixel_index2 <= 5122)) || ((pixel_index2 >= 5125) && (pixel_index2 <= 5129)) || ((pixel_index2 >= 5131) && (pixel_index2 <= 5132)) || ((pixel_index2 >= 5137) && (pixel_index2 <= 5139)) || ((pixel_index2 >= 5149) && (pixel_index2 <= 5150)) || ((pixel_index2 >= 5155) && (pixel_index2 <= 5159)) || ((pixel_index2 >= 5161) && (pixel_index2 <= 5163)) || ((pixel_index2 >= 5166) && (pixel_index2 <= 5168)) || ((pixel_index2 >= 5170) && (pixel_index2 <= 5172)) || ((pixel_index2 >= 5196) && (pixel_index2 <= 5197)) || ((pixel_index2 >= 5201) && (pixel_index2 <= 5202)) || ((pixel_index2 >= 5204) && (pixel_index2 <= 5205)) || ((pixel_index2 >= 5210) && (pixel_index2 <= 5211)) || ((pixel_index2 >= 5217) && (pixel_index2 <= 5218)) || ((pixel_index2 >= 5222) && (pixel_index2 <= 5225)) || ((pixel_index2 >= 5227) && (pixel_index2 <= 5228)) || ((pixel_index2 >= 5234) && (pixel_index2 <= 5235)) || ((pixel_index2 >= 5245) && (pixel_index2 <= 5246)) || ((pixel_index2 >= 5252) && (pixel_index2 <= 5255)) || ((pixel_index2 >= 5257) && (pixel_index2 <= 5258)) || ((pixel_index2 >= 5263) && (pixel_index2 <= 5264)) || ((pixel_index2 >= 5266) && (pixel_index2 <= 5267)) || ((pixel_index2 >= 5292) && (pixel_index2 <= 5293)) || ((pixel_index2 >= 5297) && (pixel_index2 <= 5298)) || ((pixel_index2 >= 5300) && (pixel_index2 <= 5301)) || ((pixel_index2 >= 5306) && (pixel_index2 <= 5307)) || ((pixel_index2 >= 5313) && (pixel_index2 <= 5314)) || ((pixel_index2 >= 5317) && (pixel_index2 <= 5321)) || ((pixel_index2 >= 5323) && (pixel_index2 <= 5324)) || ((pixel_index2 >= 5330) && (pixel_index2 <= 5331)) || ((pixel_index2 >= 5341) && (pixel_index2 <= 5342)) || ((pixel_index2 >= 5347) && (pixel_index2 <= 5351)) || ((pixel_index2 >= 5353) && (pixel_index2 <= 5354)) || ((pixel_index2 >= 5359) && (pixel_index2 <= 5360)) || ((pixel_index2 >= 5362) && (pixel_index2 <= 5366)) || ((pixel_index2 >= 5388) && (pixel_index2 <= 5389)) || ((pixel_index2 >= 5393) && (pixel_index2 <= 5394)) || ((pixel_index2 >= 5396) && (pixel_index2 <= 5397)) || ((pixel_index2 >= 5402) && (pixel_index2 <= 5403)) || ((pixel_index2 >= 5409) && (pixel_index2 <= 5410)) || ((pixel_index2 >= 5412) && (pixel_index2 <= 5414)) || ((pixel_index2 >= 5416) && (pixel_index2 <= 5417)) || ((pixel_index2 >= 5419) && (pixel_index2 <= 5420)) || ((pixel_index2 >= 5426) && (pixel_index2 <= 5427)) || ((pixel_index2 >= 5437) && (pixel_index2 <= 5438)) || ((pixel_index2 >= 5442) && (pixel_index2 <= 5444)) || ((pixel_index2 >= 5446) && (pixel_index2 <= 5447)) || ((pixel_index2 >= 5449) && (pixel_index2 <= 5450)) || ((pixel_index2 >= 5455) && (pixel_index2 <= 5456)) || ((pixel_index2 >= 5459) && (pixel_index2 <= 5463)) || ((pixel_index2 >= 5484) && (pixel_index2 <= 5485)) || ((pixel_index2 >= 5489) && (pixel_index2 <= 5490)) || ((pixel_index2 >= 5492) && (pixel_index2 <= 5493)) || ((pixel_index2 >= 5498) && (pixel_index2 <= 5499)) || ((pixel_index2 >= 5505) && (pixel_index2 <= 5506)) || ((pixel_index2 >= 5508) && (pixel_index2 <= 5509)) || ((pixel_index2 >= 5512) && (pixel_index2 <= 5513)) || ((pixel_index2 >= 5515) && (pixel_index2 <= 5516)) || ((pixel_index2 >= 5522) && (pixel_index2 <= 5523)) || ((pixel_index2 >= 5533) && (pixel_index2 <= 5534)) || ((pixel_index2 >= 5538) && (pixel_index2 <= 5539)) || ((pixel_index2 >= 5542) && (pixel_index2 <= 5543)) || ((pixel_index2 >= 5545) && (pixel_index2 <= 5546)) || ((pixel_index2 >= 5551) && (pixel_index2 <= 5552)) || ((pixel_index2 >= 5558) && (pixel_index2 <= 5559)) || ((pixel_index2 >= 5580) && (pixel_index2 <= 5581)) || ((pixel_index2 >= 5585) && (pixel_index2 <= 5586)) || ((pixel_index2 >= 5588) && (pixel_index2 <= 5589)) || ((pixel_index2 >= 5594) && (pixel_index2 <= 5595)) || ((pixel_index2 >= 5600) && (pixel_index2 <= 5602)) || ((pixel_index2 >= 5604) && (pixel_index2 <= 5605)) || ((pixel_index2 >= 5608) && (pixel_index2 <= 5609)) || ((pixel_index2 >= 5611) && (pixel_index2 <= 5612)) || ((pixel_index2 >= 5617) && (pixel_index2 <= 5619)) || ((pixel_index2 >= 5629) && (pixel_index2 <= 5630)) || ((pixel_index2 >= 5634) && (pixel_index2 <= 5635)) || ((pixel_index2 >= 5638) && (pixel_index2 <= 5639)) || ((pixel_index2 >= 5641) && (pixel_index2 <= 5643)) || ((pixel_index2 >= 5646) && (pixel_index2 <= 5648)) || ((pixel_index2 >= 5653) && (pixel_index2 <= 5655)) || ((pixel_index2 >= 5672) && (pixel_index2 <= 5679)) || ((pixel_index2 >= 5681) && (pixel_index2 <= 5682)) || ((pixel_index2 >= 5684) && (pixel_index2 <= 5685)) || ((pixel_index2 >= 5690) && (pixel_index2 <= 5691)) || ((pixel_index2 >= 5693) && (pixel_index2 <= 5698)) || ((pixel_index2 >= 5700) && (pixel_index2 <= 5705)) || ((pixel_index2 >= 5707) && (pixel_index2 <= 5708)) || ((pixel_index2 >= 5710) && (pixel_index2 <= 5715)) || ((pixel_index2 >= 5721) && (pixel_index2 <= 5728)) || ((pixel_index2 >= 5730) && (pixel_index2 <= 5735)) || ((pixel_index2 >= 5737) && (pixel_index2 <= 5744)) || ((pixel_index2 >= 5746) && (pixel_index2 <= 5751)) || ((pixel_index2 >= 5769) && (pixel_index2 <= 5774)) || pixel_index2 == 5777 || pixel_index2 == 5781 || pixel_index2 == 5786 || ((pixel_index2 >= 5790) && (pixel_index2 <= 5793)) || ((pixel_index2 >= 5797) && (pixel_index2 <= 5800)) || pixel_index2 == 5803 || ((pixel_index2 >= 5807) && (pixel_index2 <= 5810)) || ((pixel_index2 >= 5818) && (pixel_index2 <= 5823)) || ((pixel_index2 >= 5827) && (pixel_index2 <= 5830)) || ((pixel_index2 >= 5834) && (pixel_index2 <= 5839)) || (pixel_index2 >= 5843) && (pixel_index2 <= 5846)) oled_data2 = 16'b1111010100010100;
                    else oled_data2 = 0;
                end
                4: begin
                    if (pixel_index2 == 97 || pixel_index2 == 99 || pixel_index2 == 101 || ((pixel_index2 >= 103) && (pixel_index2 <= 104)) || ((pixel_index2 >= 106) && (pixel_index2 <= 109)) || pixel_index2 == 111 || ((pixel_index2 >= 113) && (pixel_index2 <= 114)) || ((pixel_index2 >= 118) && (pixel_index2 <= 120)) || ((pixel_index2 >= 129) && (pixel_index2 <= 165)) || pixel_index2 == 195 || pixel_index2 == 197 || ((pixel_index2 >= 199) && (pixel_index2 <= 200)) || pixel_index2 == 202 || ((pixel_index2 >= 204) && (pixel_index2 <= 205)) || pixel_index2 == 207 || ((pixel_index2 >= 209) && (pixel_index2 <= 210)) || pixel_index2 == 213 || pixel_index2 == 225 || pixel_index2 == 261 || pixel_index2 == 289 || ((pixel_index2 >= 291) && (pixel_index2 <= 296)) || pixel_index2 == 298 || ((pixel_index2 >= 300) && (pixel_index2 <= 301)) || pixel_index2 == 303 || ((pixel_index2 >= 305) && (pixel_index2 <= 306)) || ((pixel_index2 >= 310) && (pixel_index2 <= 312)) || pixel_index2 == 321 || pixel_index2 == 357 || pixel_index2 == 385 || ((pixel_index2 >= 387) && (pixel_index2 <= 392)) || pixel_index2 == 394 || ((pixel_index2 >= 396) && (pixel_index2 <= 397)) || ((pixel_index2 >= 399) && (pixel_index2 <= 402)) || pixel_index2 == 408 || pixel_index2 == 417 || pixel_index2 == 453 || ((pixel_index2 >= 501) && (pixel_index2 <= 504)) || pixel_index2 == 513 || pixel_index2 == 549 || pixel_index2 == 609 || pixel_index2 == 645 || ((pixel_index2 >= 674) && (pixel_index2 <= 675)) || ((pixel_index2 >= 678) && (pixel_index2 <= 681)) || ((pixel_index2 >= 685) && (pixel_index2 <= 686)) || pixel_index2 == 688 || ((pixel_index2 >= 690) && (pixel_index2 <= 691)) || ((pixel_index2 >= 693) && (pixel_index2 <= 696)) || pixel_index2 == 698 || pixel_index2 == 705 || pixel_index2 == 741 || ((pixel_index2 >= 770) && (pixel_index2 <= 771)) || pixel_index2 == 774 || ((pixel_index2 >= 776) && (pixel_index2 <= 777)) || ((pixel_index2 >= 779) && (pixel_index2 <= 782)) || pixel_index2 == 784 || ((pixel_index2 >= 786) && (pixel_index2 <= 787)) || ((pixel_index2 >= 790) && (pixel_index2 <= 791)) || ((pixel_index2 >= 801) && (pixel_index2 <= 837)) || ((pixel_index2 >= 866) && (pixel_index2 <= 867)) || pixel_index2 == 870 || ((pixel_index2 >= 872) && (pixel_index2 <= 873)) || pixel_index2 == 875 || ((pixel_index2 >= 877) && (pixel_index2 <= 878)) || pixel_index2 == 880 || ((pixel_index2 >= 882) && (pixel_index2 <= 883)) || ((pixel_index2 >= 886) && (pixel_index2 <= 887)) || ((pixel_index2 >= 961) && (pixel_index2 <= 964)) || pixel_index2 == 966 || ((pixel_index2 >= 968) && (pixel_index2 <= 969)) || ((pixel_index2 >= 971) && (pixel_index2 <= 974)) || ((pixel_index2 >= 976) && (pixel_index2 <= 979)) || ((pixel_index2 >= 981) && (pixel_index2 <= 984)) || pixel_index2 == 986) oled_data2 = 16'b1111001010010100;
                    else if (((pixel_index2 >= 124) && (pixel_index2 <= 128)) || ((pixel_index2 >= 166) && (pixel_index2 <= 190)) || ((pixel_index2 >= 220) && (pixel_index2 <= 221)) || pixel_index2 == 229 || pixel_index2 == 233 || pixel_index2 == 237 || pixel_index2 == 241 || pixel_index2 == 245 || pixel_index2 == 249 || pixel_index2 == 253 || pixel_index2 == 257 || pixel_index2 == 265 || pixel_index2 == 269 || pixel_index2 == 273 || pixel_index2 == 277 || pixel_index2 == 281 || ((pixel_index2 >= 285) && (pixel_index2 <= 286)) || ((pixel_index2 >= 316) && (pixel_index2 <= 317)) || pixel_index2 == 325 || pixel_index2 == 329 || pixel_index2 == 333 || pixel_index2 == 337 || pixel_index2 == 341 || pixel_index2 == 345 || pixel_index2 == 349 || pixel_index2 == 353 || pixel_index2 == 361 || pixel_index2 == 365 || pixel_index2 == 369 || pixel_index2 == 373 || pixel_index2 == 377 || ((pixel_index2 >= 381) && (pixel_index2 <= 382)) || ((pixel_index2 >= 412) && (pixel_index2 <= 413)) || pixel_index2 == 421 || pixel_index2 == 425 || pixel_index2 == 429 || pixel_index2 == 433 || pixel_index2 == 437 || pixel_index2 == 441 || pixel_index2 == 445 || pixel_index2 == 449 || pixel_index2 == 457 || pixel_index2 == 461 || pixel_index2 == 465 || pixel_index2 == 469 || pixel_index2 == 473 || ((pixel_index2 >= 477) && (pixel_index2 <= 478)) || ((pixel_index2 >= 508) && (pixel_index2 <= 509)) || pixel_index2 == 517 || pixel_index2 == 521 || pixel_index2 == 525 || pixel_index2 == 529 || pixel_index2 == 533 || pixel_index2 == 537 || pixel_index2 == 541 || pixel_index2 == 545 || pixel_index2 == 553 || pixel_index2 == 557 || pixel_index2 == 561 || pixel_index2 == 565 || pixel_index2 == 569 || ((pixel_index2 >= 573) && (pixel_index2 <= 574)) || ((pixel_index2 >= 604) && (pixel_index2 <= 605)) || pixel_index2 == 613 || pixel_index2 == 617 || pixel_index2 == 621 || pixel_index2 == 625 || pixel_index2 == 629 || pixel_index2 == 633 || pixel_index2 == 637 || pixel_index2 == 641 || pixel_index2 == 649 || pixel_index2 == 653 || pixel_index2 == 657 || pixel_index2 == 661 || pixel_index2 == 665 || ((pixel_index2 >= 669) && (pixel_index2 <= 670)) || ((pixel_index2 >= 700) && (pixel_index2 <= 701)) || pixel_index2 == 709 || pixel_index2 == 713 || pixel_index2 == 717 || pixel_index2 == 721 || pixel_index2 == 725 || pixel_index2 == 729 || pixel_index2 == 733 || pixel_index2 == 737 || pixel_index2 == 745 || pixel_index2 == 749 || pixel_index2 == 753 || pixel_index2 == 757 || pixel_index2 == 761 || ((pixel_index2 >= 765) && (pixel_index2 <= 766)) || ((pixel_index2 >= 796) && (pixel_index2 <= 800)) || ((pixel_index2 >= 838) && (pixel_index2 <= 862)) || ((pixel_index2 >= 892) && (pixel_index2 <= 894)) || ((pixel_index2 >= 897) && (pixel_index2 <= 898)) || ((pixel_index2 >= 901) && (pixel_index2 <= 902)) || ((pixel_index2 >= 905) && (pixel_index2 <= 906)) || ((pixel_index2 >= 909) && (pixel_index2 <= 910)) || ((pixel_index2 >= 913) && (pixel_index2 <= 914)) || ((pixel_index2 >= 917) && (pixel_index2 <= 918)) || ((pixel_index2 >= 921) && (pixel_index2 <= 922)) || ((pixel_index2 >= 925) && (pixel_index2 <= 926)) || ((pixel_index2 >= 929) && (pixel_index2 <= 930)) || ((pixel_index2 >= 933) && (pixel_index2 <= 934)) || ((pixel_index2 >= 937) && (pixel_index2 <= 938)) || ((pixel_index2 >= 941) && (pixel_index2 <= 942)) || ((pixel_index2 >= 945) && (pixel_index2 <= 946)) || ((pixel_index2 >= 949) && (pixel_index2 <= 950)) || ((pixel_index2 >= 953) && (pixel_index2 <= 954)) || ((pixel_index2 >= 957) && (pixel_index2 <= 958)) || ((pixel_index2 >= 988) && (pixel_index2 <= 1054)) || ((pixel_index2 >= 1084) && (pixel_index2 <= 1085)) || ((pixel_index2 >= 1087) && (pixel_index2 <= 1089)) || ((pixel_index2 >= 1091) && (pixel_index2 <= 1093)) || ((pixel_index2 >= 1095) && (pixel_index2 <= 1097)) || ((pixel_index2 >= 1099) && (pixel_index2 <= 1101)) || ((pixel_index2 >= 1103) && (pixel_index2 <= 1105)) || ((pixel_index2 >= 1107) && (pixel_index2 <= 1109)) || ((pixel_index2 >= 1111) && (pixel_index2 <= 1113)) || ((pixel_index2 >= 1115) && (pixel_index2 <= 1117)) || ((pixel_index2 >= 1119) && (pixel_index2 <= 1121)) || ((pixel_index2 >= 1123) && (pixel_index2 <= 1125)) || ((pixel_index2 >= 1127) && (pixel_index2 <= 1129)) || ((pixel_index2 >= 1131) && (pixel_index2 <= 1133)) || ((pixel_index2 >= 1135) && (pixel_index2 <= 1137)) || ((pixel_index2 >= 1139) && (pixel_index2 <= 1141)) || ((pixel_index2 >= 1143) && (pixel_index2 <= 1145)) || ((pixel_index2 >= 1147) && (pixel_index2 <= 1150)) || ((pixel_index2 >= 1182) && (pixel_index2 <= 1219)) || ((pixel_index2 >= 1240) && (pixel_index2 <= 1244)) || ((pixel_index2 >= 1278) && (pixel_index2 <= 1280)) || ((pixel_index2 >= 1283) && (pixel_index2 <= 1286)) || ((pixel_index2 >= 1290) && (pixel_index2 <= 1291)) || ((pixel_index2 >= 1293) && (pixel_index2 <= 1294)) || ((pixel_index2 >= 1314) && (pixel_index2 <= 1315)) || ((pixel_index2 >= 1336) && (pixel_index2 <= 1340)) || ((pixel_index2 >= 1374) && (pixel_index2 <= 1376)) || ((pixel_index2 >= 1378) && (pixel_index2 <= 1382)) || ((pixel_index2 >= 1386) && (pixel_index2 <= 1390)) || ((pixel_index2 >= 1410) && (pixel_index2 <= 1411)) || ((pixel_index2 >= 1432) && (pixel_index2 <= 1436)) || ((pixel_index2 >= 1470) && (pixel_index2 <= 1478)) || ((pixel_index2 >= 1482) && (pixel_index2 <= 1486)) || ((pixel_index2 >= 1506) && (pixel_index2 <= 1507)) || ((pixel_index2 >= 1528) && (pixel_index2 <= 1532)) || ((pixel_index2 >= 1566) && (pixel_index2 <= 1577)) || ((pixel_index2 >= 1583) && (pixel_index2 <= 1603)) || ((pixel_index2 >= 1624) && (pixel_index2 <= 1628)) || ((pixel_index2 >= 1662) && (pixel_index2 <= 1666)) || pixel_index2 == 1670 || ((pixel_index2 >= 1679) && (pixel_index2 <= 1696)) || ((pixel_index2 >= 1698) && (pixel_index2 <= 1699)) || ((pixel_index2 >= 1720) && (pixel_index2 <= 1724)) || ((pixel_index2 >= 1758) && (pixel_index2 <= 1762)) || pixel_index2 == 1766 || pixel_index2 == 1775 || ((pixel_index2 >= 1777) && (pixel_index2 <= 1789)) || pixel_index2 == 1792 || ((pixel_index2 >= 1794) && (pixel_index2 <= 1795)) || pixel_index2 == 1816 || ((pixel_index2 >= 1818) && (pixel_index2 <= 1820)) || ((pixel_index2 >= 1854) && (pixel_index2 <= 1858)) || pixel_index2 == 1862 || ((pixel_index2 >= 1872) && (pixel_index2 <= 1878)) || ((pixel_index2 >= 1882) && (pixel_index2 <= 1888)) || ((pixel_index2 >= 1892) && (pixel_index2 <= 1913)) || ((pixel_index2 >= 1915) && (pixel_index2 <= 1916)) || ((pixel_index2 >= 1948) && (pixel_index2 <= 1961)) || ((pixel_index2 >= 1967) && (pixel_index2 <= 1973)) || pixel_index2 == 1988 || pixel_index2 == 1991 || ((pixel_index2 >= 1993) && (pixel_index2 <= 1994)) || pixel_index2 == 1996 || ((pixel_index2 >= 2000) && (pixel_index2 <= 2001)) || pixel_index2 == 2008 || ((pixel_index2 >= 2011) && (pixel_index2 <= 2014)) || ((pixel_index2 >= 2044) && (pixel_index2 <= 2046)) || ((pixel_index2 >= 2048) && (pixel_index2 <= 2054)) || ((pixel_index2 >= 2058) && (pixel_index2 <= 2069)) || ((pixel_index2 >= 2084) && (pixel_index2 <= 2085)) || pixel_index2 == 2089 || ((pixel_index2 >= 2091) && (pixel_index2 <= 2093)) || ((pixel_index2 >= 2095) && (pixel_index2 <= 2096)) || ((pixel_index2 >= 2104) && (pixel_index2 <= 2105)) || ((pixel_index2 >= 2107) && (pixel_index2 <= 2110)) || pixel_index2 == 2140 || pixel_index2 == 2142 || ((pixel_index2 >= 2144) && (pixel_index2 <= 2150)) || pixel_index2 == 2154 || ((pixel_index2 >= 2157) && (pixel_index2 <= 2168)) || pixel_index2 == 2178 || ((pixel_index2 >= 2180) && (pixel_index2 <= 2184)) || pixel_index2 == 2188 || ((pixel_index2 >= 2190) && (pixel_index2 <= 2192)) || ((pixel_index2 >= 2195) && (pixel_index2 <= 2197)) || ((pixel_index2 >= 2200) && (pixel_index2 <= 2206)) || ((pixel_index2 >= 2236) && (pixel_index2 <= 2238)) || ((pixel_index2 >= 2245) && (pixel_index2 <= 2246)) || pixel_index2 == 2250 || ((pixel_index2 >= 2252) && (pixel_index2 <= 2264)) || ((pixel_index2 >= 2274) && (pixel_index2 <= 2288)) || ((pixel_index2 >= 2291) && (pixel_index2 <= 2293)) || ((pixel_index2 >= 2296) && (pixel_index2 <= 2302)) || ((pixel_index2 >= 2332) && (pixel_index2 <= 2334)) || ((pixel_index2 >= 2341) && (pixel_index2 <= 2355)) || ((pixel_index2 >= 2374) && (pixel_index2 <= 2384)) || ((pixel_index2 >= 2392) && (pixel_index2 <= 2398)) || ((pixel_index2 >= 2428) && (pixel_index2 <= 2437)) || ((pixel_index2 >= 2443) && (pixel_index2 <= 2451)) || ((pixel_index2 >= 2470) && (pixel_index2 <= 2480)) || ((pixel_index2 >= 2487) && (pixel_index2 <= 2494)) || ((pixel_index2 >= 2526) && (pixel_index2 <= 2532)) || ((pixel_index2 >= 2540) && (pixel_index2 <= 2547)) || pixel_index2 == 2566 || ((pixel_index2 >= 2580) && (pixel_index2 <= 2588)) || ((pixel_index2 >= 2622) && (pixel_index2 <= 2626)) || pixel_index2 == 2636 || ((pixel_index2 >= 2639) && (pixel_index2 <= 2644)) || ((pixel_index2 >= 2647) && (pixel_index2 <= 2648)) || pixel_index2 == 2659 || ((pixel_index2 >= 2661) && (pixel_index2 <= 2662)) || ((pixel_index2 >= 2676) && (pixel_index2 <= 2684)) || ((pixel_index2 >= 2718) && (pixel_index2 <= 2721)) || pixel_index2 == 2732 || ((pixel_index2 >= 2735) && (pixel_index2 <= 2742)) || ((pixel_index2 >= 2756) && (pixel_index2 <= 2758)) || ((pixel_index2 >= 2772) && (pixel_index2 <= 2780)) || ((pixel_index2 >= 2814) && (pixel_index2 <= 2817)) || pixel_index2 == 2828 || ((pixel_index2 >= 2831) && (pixel_index2 <= 2838)) || ((pixel_index2 >= 2842) && (pixel_index2 <= 2848)) || ((pixel_index2 >= 2852) && (pixel_index2 <= 2859)) || ((pixel_index2 >= 2866) && (pixel_index2 <= 2876)) || ((pixel_index2 >= 2910) && (pixel_index2 <= 2913)) || pixel_index2 == 2924 || ((pixel_index2 >= 2927) && (pixel_index2 <= 2935)) || ((pixel_index2 >= 2938) && (pixel_index2 <= 2944)) || ((pixel_index2 >= 2947) && (pixel_index2 <= 2955)) || pixel_index2 == 2962 || ((pixel_index2 >= 2964) && (pixel_index2 <= 2972)) || ((pixel_index2 >= 3006) && (pixel_index2 <= 3013)) || ((pixel_index2 >= 3019) && (pixel_index2 <= 3021)) || ((pixel_index2 >= 3023) && (pixel_index2 <= 3032)) || ((pixel_index2 >= 3042) && (pixel_index2 <= 3051)) || ((pixel_index2 >= 3058) && (pixel_index2 <= 3060)) || pixel_index2 == 3063 || ((pixel_index2 >= 3065) && (pixel_index2 <= 3068)) || ((pixel_index2 >= 3102) && (pixel_index2 <= 3104)) || pixel_index2 == 3107 || ((pixel_index2 >= 3117) && (pixel_index2 <= 3123)) || ((pixel_index2 >= 3143) && (pixel_index2 <= 3147)) || ((pixel_index2 >= 3154) && (pixel_index2 <= 3155)) || pixel_index2 == 3159 || ((pixel_index2 >= 3161) && (pixel_index2 <= 3164)) || ((pixel_index2 >= 3198) && (pixel_index2 <= 3200)) || ((pixel_index2 >= 3202) && (pixel_index2 <= 3203)) || ((pixel_index2 >= 3213) && (pixel_index2 <= 3216)) || ((pixel_index2 >= 3218) && (pixel_index2 <= 3219)) || ((pixel_index2 >= 3239) && (pixel_index2 <= 3243)) || ((pixel_index2 >= 3250) && (pixel_index2 <= 3251)) || ((pixel_index2 >= 3255) && (pixel_index2 <= 3260)) || ((pixel_index2 >= 3292) && (pixel_index2 <= 3299)) || ((pixel_index2 >= 3309) && (pixel_index2 <= 3312)) || ((pixel_index2 >= 3314) && (pixel_index2 <= 3315)) || ((pixel_index2 >= 3335) && (pixel_index2 <= 3337)) || pixel_index2 == 3339 || ((pixel_index2 >= 3346) && (pixel_index2 <= 3347)) || ((pixel_index2 >= 3351) && (pixel_index2 <= 3352)) || ((pixel_index2 >= 3354) && (pixel_index2 <= 3358)) || ((pixel_index2 >= 3388) && (pixel_index2 <= 3393)) || pixel_index2 == 3395 || ((pixel_index2 >= 3405) && (pixel_index2 <= 3407)) || ((pixel_index2 >= 3409) && (pixel_index2 <= 3411)) || ((pixel_index2 >= 3431) && (pixel_index2 <= 3432)) || ((pixel_index2 >= 3434) && (pixel_index2 <= 3435)) || ((pixel_index2 >= 3438) && (pixel_index2 <= 3443)) || ((pixel_index2 >= 3447) && (pixel_index2 <= 3448)) || ((pixel_index2 >= 3450) && (pixel_index2 <= 3454)) || ((pixel_index2 >= 3484) && (pixel_index2 <= 3487)) || pixel_index2 == 3489 || pixel_index2 == 3491 || ((pixel_index2 >= 3501) && (pixel_index2 <= 3502)) || ((pixel_index2 >= 3505) && (pixel_index2 <= 3507)) || ((pixel_index2 >= 3527) && (pixel_index2 <= 3531)) || ((pixel_index2 >= 3538) && (pixel_index2 <= 3539)) || ((pixel_index2 >= 3543) && (pixel_index2 <= 3544)) || ((pixel_index2 >= 3546) && (pixel_index2 <= 3550)) || ((pixel_index2 >= 3580) && (pixel_index2 <= 3587)) || ((pixel_index2 >= 3597) && (pixel_index2 <= 3603)) || ((pixel_index2 >= 3623) && (pixel_index2 <= 3628)) || ((pixel_index2 >= 3633) && (pixel_index2 <= 3635)) || ((pixel_index2 >= 3639) && (pixel_index2 <= 3646)) || ((pixel_index2 >= 4620) && (pixel_index2 <= 4692)) || ((pixel_index2 >= 4707) && (pixel_index2 <= 4796)) || ((pixel_index2 >= 4803) && (pixel_index2 <= 4812)) || ((pixel_index2 >= 4814) && (pixel_index2 <= 4817)) || ((pixel_index2 >= 4819) && (pixel_index2 <= 4820)) || ((pixel_index2 >= 4827) && (pixel_index2 <= 4829)) || ((pixel_index2 >= 4834) && (pixel_index2 <= 4835)) || ((pixel_index2 >= 4838) && (pixel_index2 <= 4839)) || ((pixel_index2 >= 4841) && (pixel_index2 <= 4843)) || ((pixel_index2 >= 4845) && (pixel_index2 <= 4846)) || ((pixel_index2 >= 4851) && (pixel_index2 <= 4861)) || ((pixel_index2 >= 4863) && (pixel_index2 <= 4865)) || ((pixel_index2 >= 4868) && (pixel_index2 <= 4869)) || ((pixel_index2 >= 4871) && (pixel_index2 <= 4873)) || ((pixel_index2 >= 4880) && (pixel_index2 <= 4882)) || ((pixel_index2 >= 4887) && (pixel_index2 <= 4892)) || ((pixel_index2 >= 4899) && (pixel_index2 <= 4907)) || ((pixel_index2 >= 4910) && (pixel_index2 <= 4912)) || pixel_index2 == 4915 || pixel_index2 == 4924 || pixel_index2 == 4931 || pixel_index2 == 4935 || pixel_index2 == 4938 || pixel_index2 == 4941 || ((pixel_index2 >= 4948) && (pixel_index2 <= 4956)) || ((pixel_index2 >= 4959) && (pixel_index2 <= 4961)) || pixel_index2 == 4965 || pixel_index2 == 4968 || pixel_index2 == 4977 || ((pixel_index2 >= 4984) && (pixel_index2 <= 4988)) || ((pixel_index2 >= 4994) && (pixel_index2 <= 5003)) || ((pixel_index2 >= 5006) && (pixel_index2 <= 5008)) || pixel_index2 == 5011 || pixel_index2 == 5020 || pixel_index2 == 5027 || pixel_index2 == 5034 || pixel_index2 == 5037 || ((pixel_index2 >= 5044) && (pixel_index2 <= 5052)) || ((pixel_index2 >= 5055) && (pixel_index2 <= 5057)) || pixel_index2 == 5064 || pixel_index2 == 5073 || ((pixel_index2 >= 5080) && (pixel_index2 <= 5085)) || ((pixel_index2 >= 5090) && (pixel_index2 <= 5099)) || ((pixel_index2 >= 5102) && (pixel_index2 <= 5104)) || pixel_index2 == 5107 || ((pixel_index2 >= 5111) && (pixel_index2 <= 5112)) || ((pixel_index2 >= 5116) && (pixel_index2 <= 5119)) || ((pixel_index2 >= 5123) && (pixel_index2 <= 5124)) || pixel_index2 == 5130 || ((pixel_index2 >= 5133) && (pixel_index2 <= 5136)) || ((pixel_index2 >= 5140) && (pixel_index2 <= 5148)) || ((pixel_index2 >= 5151) && (pixel_index2 <= 5154)) || pixel_index2 == 5160 || ((pixel_index2 >= 5164) && (pixel_index2 <= 5165)) || pixel_index2 == 5169 || ((pixel_index2 >= 5173) && (pixel_index2 <= 5181)) || ((pixel_index2 >= 5186) && (pixel_index2 <= 5195)) || ((pixel_index2 >= 5198) && (pixel_index2 <= 5200)) || pixel_index2 == 5203 || ((pixel_index2 >= 5206) && (pixel_index2 <= 5209)) || ((pixel_index2 >= 5212) && (pixel_index2 <= 5216)) || ((pixel_index2 >= 5219) && (pixel_index2 <= 5220)) || pixel_index2 == 5226 || ((pixel_index2 >= 5229) && (pixel_index2 <= 5233)) || ((pixel_index2 >= 5236) && (pixel_index2 <= 5244)) || ((pixel_index2 >= 5247) && (pixel_index2 <= 5250)) || pixel_index2 == 5256 || ((pixel_index2 >= 5259) && (pixel_index2 <= 5262)) || pixel_index2 == 5265 || ((pixel_index2 >= 5271) && (pixel_index2 <= 5277)) || ((pixel_index2 >= 5282) && (pixel_index2 <= 5291)) || ((pixel_index2 >= 5294) && (pixel_index2 <= 5296)) || pixel_index2 == 5299 || ((pixel_index2 >= 5302) && (pixel_index2 <= 5305)) || ((pixel_index2 >= 5308) && (pixel_index2 <= 5312)) || pixel_index2 == 5315 || pixel_index2 == 5322 || ((pixel_index2 >= 5325) && (pixel_index2 <= 5329)) || ((pixel_index2 >= 5332) && (pixel_index2 <= 5340)) || ((pixel_index2 >= 5343) && (pixel_index2 <= 5345)) || pixel_index2 == 5352 || ((pixel_index2 >= 5355) && (pixel_index2 <= 5358)) || pixel_index2 == 5361 || ((pixel_index2 >= 5368) && (pixel_index2 <= 5373)) || ((pixel_index2 >= 5378) && (pixel_index2 <= 5387)) || ((pixel_index2 >= 5390) && (pixel_index2 <= 5392)) || pixel_index2 == 5395 || ((pixel_index2 >= 5398) && (pixel_index2 <= 5401)) || ((pixel_index2 >= 5404) && (pixel_index2 <= 5408)) || pixel_index2 == 5411 || pixel_index2 == 5415 || pixel_index2 == 5418 || ((pixel_index2 >= 5421) && (pixel_index2 <= 5425)) || ((pixel_index2 >= 5428) && (pixel_index2 <= 5436)) || ((pixel_index2 >= 5439) && (pixel_index2 <= 5441)) || pixel_index2 == 5445 || pixel_index2 == 5448 || ((pixel_index2 >= 5451) && (pixel_index2 <= 5454)) || ((pixel_index2 >= 5457) && (pixel_index2 <= 5458)) || ((pixel_index2 >= 5464) && (pixel_index2 <= 5469)) || ((pixel_index2 >= 5474) && (pixel_index2 <= 5483)) || ((pixel_index2 >= 5486) && (pixel_index2 <= 5488)) || pixel_index2 == 5491 || ((pixel_index2 >= 5494) && (pixel_index2 <= 5497)) || ((pixel_index2 >= 5500) && (pixel_index2 <= 5503)) || pixel_index2 == 5507 || ((pixel_index2 >= 5510) && (pixel_index2 <= 5511)) || pixel_index2 == 5514 || ((pixel_index2 >= 5517) && (pixel_index2 <= 5520)) || ((pixel_index2 >= 5524) && (pixel_index2 <= 5532)) || ((pixel_index2 >= 5535) && (pixel_index2 <= 5537)) || ((pixel_index2 >= 5540) && (pixel_index2 <= 5541)) || pixel_index2 == 5544 || ((pixel_index2 >= 5548) && (pixel_index2 <= 5549)) || ((pixel_index2 >= 5553) && (pixel_index2 <= 5556)) || ((pixel_index2 >= 5560) && (pixel_index2 <= 5565)) || ((pixel_index2 >= 5570) && (pixel_index2 <= 5575)) || pixel_index2 == 5584 || pixel_index2 == 5587 || ((pixel_index2 >= 5590) && (pixel_index2 <= 5593)) || pixel_index2 == 5596 || pixel_index2 == 5603 || pixel_index2 == 5610 || pixel_index2 == 5613 || ((pixel_index2 >= 5620) && (pixel_index2 <= 5624)) || pixel_index2 == 5633 || pixel_index2 == 5640 || pixel_index2 == 5649 || ((pixel_index2 >= 5656) && (pixel_index2 <= 5661)) || ((pixel_index2 >= 5667) && (pixel_index2 <= 5671)) || pixel_index2 == 5680 || pixel_index2 == 5683 || ((pixel_index2 >= 5686) && (pixel_index2 <= 5689)) || pixel_index2 == 5692 || pixel_index2 == 5699 || pixel_index2 == 5706 || pixel_index2 == 5709 || ((pixel_index2 >= 5716) && (pixel_index2 <= 5720)) || pixel_index2 == 5729 || pixel_index2 == 5736 || pixel_index2 == 5745 || ((pixel_index2 >= 5752) && (pixel_index2 <= 5756)) || ((pixel_index2 >= 5763) && (pixel_index2 <= 5768)) || ((pixel_index2 >= 5775) && (pixel_index2 <= 5776)) || ((pixel_index2 >= 5778) && (pixel_index2 <= 5780)) || ((pixel_index2 >= 5782) && (pixel_index2 <= 5785)) || ((pixel_index2 >= 5787) && (pixel_index2 <= 5789)) || ((pixel_index2 >= 5794) && (pixel_index2 <= 5796)) || ((pixel_index2 >= 5801) && (pixel_index2 <= 5802)) || ((pixel_index2 >= 5804) && (pixel_index2 <= 5806)) || ((pixel_index2 >= 5811) && (pixel_index2 <= 5817)) || ((pixel_index2 >= 5824) && (pixel_index2 <= 5826)) || ((pixel_index2 >= 5831) && (pixel_index2 <= 5833)) || ((pixel_index2 >= 5840) && (pixel_index2 <= 5842)) || ((pixel_index2 >= 5847) && (pixel_index2 <= 5852)) || (pixel_index2 >= 5868) && (pixel_index2 <= 5940)) oled_data2 = 16'b0000000000001010;
                    else if (pixel_index2 == 339 || pixel_index2 == 343 || pixel_index2 == 347 || pixel_index2 == 351 || pixel_index2 == 355 || pixel_index2 == 435 || pixel_index2 == 439 || pixel_index2 == 443 || pixel_index2 == 447 || pixel_index2 == 451 || pixel_index2 == 3253 || pixel_index2 == 3349) oled_data2 = 16'b0000010100000000;
                    else if (pixel_index2 == 511 || pixel_index2 == 515 || pixel_index2 == 519 || pixel_index2 == 523 || pixel_index2 == 527 || pixel_index2 == 551 || pixel_index2 == 555 || pixel_index2 == 559 || pixel_index2 == 563 || pixel_index2 == 567 || pixel_index2 == 571 || pixel_index2 == 607 || pixel_index2 == 611 || pixel_index2 == 615 || pixel_index2 == 619 || pixel_index2 == 623 || pixel_index2 == 647 || pixel_index2 == 651 || pixel_index2 == 655 || pixel_index2 == 659 || pixel_index2 == 663 || pixel_index2 == 667 || pixel_index2 == 3488) oled_data2 = 16'b1010000000000000;
                    else if (((pixel_index2 >= 895) && (pixel_index2 <= 896)) || ((pixel_index2 >= 899) && (pixel_index2 <= 900)) || ((pixel_index2 >= 903) && (pixel_index2 <= 904)) || ((pixel_index2 >= 907) && (pixel_index2 <= 908)) || ((pixel_index2 >= 911) && (pixel_index2 <= 912)) || ((pixel_index2 >= 915) && (pixel_index2 <= 916)) || ((pixel_index2 >= 919) && (pixel_index2 <= 920)) || ((pixel_index2 >= 923) && (pixel_index2 <= 924)) || ((pixel_index2 >= 927) && (pixel_index2 <= 928)) || ((pixel_index2 >= 931) && (pixel_index2 <= 932)) || ((pixel_index2 >= 935) && (pixel_index2 <= 936)) || ((pixel_index2 >= 939) && (pixel_index2 <= 940)) || ((pixel_index2 >= 943) && (pixel_index2 <= 944)) || ((pixel_index2 >= 947) && (pixel_index2 <= 948)) || ((pixel_index2 >= 951) && (pixel_index2 <= 952)) || ((pixel_index2 >= 955) && (pixel_index2 <= 956)) || pixel_index2 == 1155 || ((pixel_index2 >= 1159) && (pixel_index2 <= 1161)) || pixel_index2 == 1163 || ((pixel_index2 >= 1165) && (pixel_index2 <= 1166)) || pixel_index2 == 1168 || ((pixel_index2 >= 1170) && (pixel_index2 <= 1171)) || pixel_index2 == 1173 || ((pixel_index2 >= 1175) && (pixel_index2 <= 1176)) || pixel_index2 == 1254 || ((pixel_index2 >= 1256) && (pixel_index2 <= 1257)) || pixel_index2 == 1259 || ((pixel_index2 >= 1261) && (pixel_index2 <= 1262)) || ((pixel_index2 >= 1264) && (pixel_index2 <= 1267)) || ((pixel_index2 >= 1270) && (pixel_index2 <= 1272)) || pixel_index2 == 1350 || ((pixel_index2 >= 1352) && (pixel_index2 <= 1353)) || pixel_index2 == 1355 || ((pixel_index2 >= 1357) && (pixel_index2 <= 1358)) || pixel_index2 == 1360 || ((pixel_index2 >= 1362) && (pixel_index2 <= 1363)) || pixel_index2 == 1365 || ((pixel_index2 >= 1367) && (pixel_index2 <= 1368)) || ((pixel_index2 >= 1447) && (pixel_index2 <= 1449)) || ((pixel_index2 >= 1451) && (pixel_index2 <= 1454)) || ((pixel_index2 >= 1456) && (pixel_index2 <= 1459)) || ((pixel_index2 >= 1461) && (pixel_index2 <= 1464)) || ((pixel_index2 >= 1637) && (pixel_index2 <= 1638)) || ((pixel_index2 >= 1641) && (pixel_index2 <= 1644)) || ((pixel_index2 >= 1646) && (pixel_index2 <= 1649)) || ((pixel_index2 >= 1652) && (pixel_index2 <= 1654)) || pixel_index2 == 1732 || pixel_index2 == 1735 || pixel_index2 == 1740 || pixel_index2 == 1745 || pixel_index2 == 1747 || pixel_index2 == 1831 || pixel_index2 == 1836 || ((pixel_index2 >= 1839) && (pixel_index2 <= 1841)) || ((pixel_index2 >= 1844) && (pixel_index2 <= 1845)) || pixel_index2 == 1924 || pixel_index2 == 1927 || pixel_index2 == 1932 || pixel_index2 == 1937 || pixel_index2 == 1942 || ((pixel_index2 >= 2021) && (pixel_index2 <= 2022)) || pixel_index2 == 2028 || ((pixel_index2 >= 2030) && (pixel_index2 <= 2033)) || ((pixel_index2 >= 2035) && (pixel_index2 <= 2037)) || pixel_index2 == 2213 || pixel_index2 == 2216 || ((pixel_index2 >= 2219) && (pixel_index2 <= 2221)) || pixel_index2 == 2223 || pixel_index2 == 2226 || ((pixel_index2 >= 2228) && (pixel_index2 <= 2230)) || pixel_index2 == 2310 || pixel_index2 == 2312 || pixel_index2 == 2314 || pixel_index2 == 2319 || pixel_index2 == 2322 || pixel_index2 == 2325 || ((pixel_index2 >= 2406) && (pixel_index2 <= 2408)) || ((pixel_index2 >= 2411) && (pixel_index2 <= 2412)) || ((pixel_index2 >= 2415) && (pixel_index2 <= 2416)) || pixel_index2 == 2418 || pixel_index2 == 2421 || pixel_index2 == 2501 || pixel_index2 == 2504 || pixel_index2 == 2509 || pixel_index2 == 2511 || ((pixel_index2 >= 2513) && (pixel_index2 <= 2514)) || pixel_index2 == 2517 || ((pixel_index2 >= 2598) && (pixel_index2 <= 2600)) || ((pixel_index2 >= 2602) && (pixel_index2 <= 2604)) || pixel_index2 == 2607 || pixel_index2 == 2610 || ((pixel_index2 >= 2612) && (pixel_index2 <= 2614)) || ((pixel_index2 >= 3133) && (pixel_index2 <= 3134)) || pixel_index2 == 3228 || pixel_index2 == 3327 || ((pixel_index2 >= 3364) && (pixel_index2 <= 3367)) || ((pixel_index2 >= 3370) && (pixel_index2 <= 3372)) || ((pixel_index2 >= 3375) && (pixel_index2 <= 3376)) || ((pixel_index2 >= 3380) && (pixel_index2 <= 3382)) || pixel_index2 == 3463 || pixel_index2 == 3465 || pixel_index2 == 3468 || pixel_index2 == 3470 || pixel_index2 == 3473 || pixel_index2 == 3475 || pixel_index2 == 3478 || pixel_index2 == 3559 || ((pixel_index2 >= 3562) && (pixel_index2 <= 3564)) || pixel_index2 == 3566 || pixel_index2 == 3569 || ((pixel_index2 >= 3572) && (pixel_index2 <= 3574)) || ((pixel_index2 >= 3630) && (pixel_index2 <= 3631)) || pixel_index2 == 3655 || pixel_index2 == 3657 || pixel_index2 == 3660 || pixel_index2 == 3662 || pixel_index2 == 3665 || pixel_index2 == 3667 || pixel_index2 == 3670 || pixel_index2 == 3751 || ((pixel_index2 >= 3754) && (pixel_index2 <= 3756)) || pixel_index2 == 3758 || pixel_index2 == 3761 || ((pixel_index2 >= 3764) && (pixel_index2 <= 3766)) || ((pixel_index2 >= 3938) && (pixel_index2 <= 3939)) || pixel_index2 == 3942 || pixel_index2 == 3945 || ((pixel_index2 >= 3947) && (pixel_index2 <= 3950)) || pixel_index2 == 3952 || ((pixel_index2 >= 3954) && (pixel_index2 <= 3955)) || ((pixel_index2 >= 3959) && (pixel_index2 <= 3962)) || ((pixel_index2 >= 3964) && (pixel_index2 <= 3967)) || ((pixel_index2 >= 3969) && (pixel_index2 <= 3972)) || ((pixel_index2 >= 3974) && (pixel_index2 <= 3977)) || pixel_index2 == 3979 || ((pixel_index2 >= 3981) && (pixel_index2 <= 3982)) || ((pixel_index2 >= 3984) && (pixel_index2 <= 3986)) || ((pixel_index2 >= 4008) && (pixel_index2 <= 4009)) || ((pixel_index2 >= 4012) && (pixel_index2 <= 4015)) || ((pixel_index2 >= 4017) && (pixel_index2 <= 4020)) || ((pixel_index2 >= 4022) && (pixel_index2 <= 4025)) || pixel_index2 == 4027 || ((pixel_index2 >= 4029) && (pixel_index2 <= 4030)) || ((pixel_index2 >= 4034) && (pixel_index2 <= 4035)) || ((pixel_index2 >= 4039) && (pixel_index2 <= 4040)) || ((pixel_index2 >= 4045) && (pixel_index2 <= 4046)) || pixel_index2 == 4048 || ((pixel_index2 >= 4050) && (pixel_index2 <= 4051)) || ((pixel_index2 >= 4057) && (pixel_index2 <= 4058)) || ((pixel_index2 >= 4060) && (pixel_index2 <= 4061)) || pixel_index2 == 4065 || ((pixel_index2 >= 4067) && (pixel_index2 <= 4068)) || pixel_index2 == 4070 || ((pixel_index2 >= 4072) && (pixel_index2 <= 4073)) || ((pixel_index2 >= 4075) && (pixel_index2 <= 4078)) || ((pixel_index2 >= 4082) && (pixel_index2 <= 4083)) || ((pixel_index2 >= 4104) && (pixel_index2 <= 4105)) || ((pixel_index2 >= 4110) && (pixel_index2 <= 4111)) || ((pixel_index2 >= 4113) && (pixel_index2 <= 4114)) || ((pixel_index2 >= 4120) && (pixel_index2 <= 4121)) || ((pixel_index2 >= 4124) && (pixel_index2 <= 4126)) || ((pixel_index2 >= 4130) && (pixel_index2 <= 4131)) || ((pixel_index2 >= 4135) && (pixel_index2 <= 4136)) || ((pixel_index2 >= 4139) && (pixel_index2 <= 4140)) || pixel_index2 == 4142 || pixel_index2 == 4144 || ((pixel_index2 >= 4146) && (pixel_index2 <= 4147)) || ((pixel_index2 >= 4151) && (pixel_index2 <= 4152)) || pixel_index2 == 4154 || ((pixel_index2 >= 4157) && (pixel_index2 <= 4159)) || pixel_index2 == 4161 || ((pixel_index2 >= 4163) && (pixel_index2 <= 4164)) || pixel_index2 == 4166 || ((pixel_index2 >= 4168) && (pixel_index2 <= 4169)) || pixel_index2 == 4171 || ((pixel_index2 >= 4173) && (pixel_index2 <= 4174)) || ((pixel_index2 >= 4178) && (pixel_index2 <= 4179)) || ((pixel_index2 >= 4200) && (pixel_index2 <= 4201)) || ((pixel_index2 >= 4204) && (pixel_index2 <= 4205)) || pixel_index2 == 4207 || ((pixel_index2 >= 4210) && (pixel_index2 <= 4212)) || ((pixel_index2 >= 4214) && (pixel_index2 <= 4215)) || pixel_index2 == 4217 || pixel_index2 == 4219 || ((pixel_index2 >= 4221) && (pixel_index2 <= 4222)) || ((pixel_index2 >= 4225) && (pixel_index2 <= 4228)) || pixel_index2 == 4230 || pixel_index2 == 4233 || ((pixel_index2 >= 4235) && (pixel_index2 <= 4238)) || ((pixel_index2 >= 4240) && (pixel_index2 <= 4243)) || ((pixel_index2 >= 4247) && (pixel_index2 <= 4250)) || ((pixel_index2 >= 4252) && (pixel_index2 <= 4254)) || ((pixel_index2 >= 4257) && (pixel_index2 <= 4260)) || ((pixel_index2 >= 4262) && (pixel_index2 <= 4265)) || pixel_index2 == 4267 || ((pixel_index2 >= 4269) && (pixel_index2 <= 4270)) || ((pixel_index2 >= 4272) && (pixel_index2 <= 4274)) || ((pixel_index2 >= 4295) && (pixel_index2 <= 4298)) || ((pixel_index2 >= 4300) && (pixel_index2 <= 4303)) || ((pixel_index2 >= 4305) && (pixel_index2 <= 4307)) || ((pixel_index2 >= 4310) && (pixel_index2 <= 4313)) || ((pixel_index2 >= 4315) && (pixel_index2 <= 4318)) || pixel_index2 == 4802 || pixel_index2 == 4893 || pixel_index2 == 5762 || pixel_index2 == 5853) oled_data2 = 16'b1111011110011110;
                    else if (pixel_index2 == 1086 || pixel_index2 == 1090 || pixel_index2 == 1094 || pixel_index2 == 1098 || pixel_index2 == 1102 || pixel_index2 == 1126 || pixel_index2 == 1130 || pixel_index2 == 1134 || pixel_index2 == 1138 || pixel_index2 == 1142 || pixel_index2 == 1146) oled_data2 = 16'b0000001010000000;
                    else if (pixel_index2 == 1106 || pixel_index2 == 1110 || pixel_index2 == 1114 || pixel_index2 == 1118 || pixel_index2 == 1122) oled_data2 = 16'b1111011110001010;
                    else if (((pixel_index2 >= 1281) && (pixel_index2 <= 1282)) || pixel_index2 == 1292 || pixel_index2 == 1295 || ((pixel_index2 >= 1297) && (pixel_index2 <= 1299)) || pixel_index2 == 1302 || ((pixel_index2 >= 1304) && (pixel_index2 <= 1305)) || pixel_index2 == 1307 || pixel_index2 == 1309 || pixel_index2 == 1311 || pixel_index2 == 1313 || pixel_index2 == 1377 || ((pixel_index2 >= 1392) && (pixel_index2 <= 1395)) || ((pixel_index2 >= 1397) && (pixel_index2 <= 1399)) || pixel_index2 == 1401 || ((pixel_index2 >= 1403) && (pixel_index2 <= 1404)) || pixel_index2 == 1406 || pixel_index2 == 1409 || ((pixel_index2 >= 1487) && (pixel_index2 <= 1488)) || pixel_index2 == 1490 || pixel_index2 == 1493 || pixel_index2 == 1495 || pixel_index2 == 1497 || ((pixel_index2 >= 1499) && (pixel_index2 <= 1500)) || ((pixel_index2 >= 1502) && (pixel_index2 <= 1503)) || pixel_index2 == 1505 || pixel_index2 == 1697 || pixel_index2 == 1776 || ((pixel_index2 >= 1790) && (pixel_index2 <= 1791)) || pixel_index2 == 1793 || pixel_index2 == 1817 || pixel_index2 == 1871 || pixel_index2 == 1914 || pixel_index2 == 1974 || ((pixel_index2 >= 1989) && (pixel_index2 <= 1990)) || pixel_index2 == 1992 || pixel_index2 == 1995 || ((pixel_index2 >= 1997) && (pixel_index2 <= 1999)) || ((pixel_index2 >= 2009) && (pixel_index2 <= 2010)) || pixel_index2 == 2047 || ((pixel_index2 >= 2070) && (pixel_index2 <= 2071)) || pixel_index2 == 2083 || ((pixel_index2 >= 2086) && (pixel_index2 <= 2088)) || pixel_index2 == 2090 || pixel_index2 == 2094 || pixel_index2 == 2106 || pixel_index2 == 2141 || pixel_index2 == 2143 || ((pixel_index2 >= 2155) && (pixel_index2 <= 2156)) || pixel_index2 == 2179 || ((pixel_index2 >= 2185) && (pixel_index2 <= 2187)) || pixel_index2 == 2189 || pixel_index2 == 2240 || pixel_index2 == 2243 || pixel_index2 == 2251 || pixel_index2 == 2336 || pixel_index2 == 2338 || pixel_index2 == 2340 || pixel_index2 == 2548 || ((pixel_index2 >= 2550) && (pixel_index2 <= 2551)) || ((pixel_index2 >= 2562) && (pixel_index2 <= 2563)) || ((pixel_index2 >= 2567) && (pixel_index2 <= 2579)) || ((pixel_index2 >= 2645) && (pixel_index2 <= 2646)) || pixel_index2 == 2658 || pixel_index2 == 2660 || ((pixel_index2 >= 2663) && (pixel_index2 <= 2675)) || ((pixel_index2 >= 2759) && (pixel_index2 <= 2771)) || ((pixel_index2 >= 2925) && (pixel_index2 <= 2926)) || pixel_index2 == 2937 || pixel_index2 == 2946 || pixel_index2 == 3022 || ((pixel_index2 >= 3105) && (pixel_index2 <= 3106)) || pixel_index2 == 3201 || pixel_index2 == 3217 || ((pixel_index2 >= 3230) && (pixel_index2 <= 3231)) || pixel_index2 == 3313 || pixel_index2 == 3324 || pixel_index2 == 3408 || ((pixel_index2 >= 3421) && (pixel_index2 <= 3422)) || ((pixel_index2 >= 3503) && (pixel_index2 <= 3504)) || ((pixel_index2 >= 3533) && (pixel_index2 <= 3536)) || pixel_index2 == 3629 || pixel_index2 == 3632) oled_data2 = 16'b1010010100010100;
                    else if (pixel_index2 == 1287 || pixel_index2 == 1289 || pixel_index2 == 1479 || pixel_index2 == 1481 || pixel_index2 == 1667 || pixel_index2 == 1669 || pixel_index2 == 1671 || pixel_index2 == 1673 || pixel_index2 == 1675 || pixel_index2 == 1677 || pixel_index2 == 1859 || pixel_index2 == 1861 || pixel_index2 == 1863 || pixel_index2 == 1865 || pixel_index2 == 1867 || pixel_index2 == 1869 || ((pixel_index2 >= 1879) && (pixel_index2 <= 1881)) || ((pixel_index2 >= 1889) && (pixel_index2 <= 1891)) || ((pixel_index2 >= 1975) && (pixel_index2 <= 1987)) || ((pixel_index2 >= 2002) && (pixel_index2 <= 2007)) || pixel_index2 == 2055 || pixel_index2 == 2057 || ((pixel_index2 >= 2072) && (pixel_index2 <= 2073)) || ((pixel_index2 >= 2081) && (pixel_index2 <= 2082)) || ((pixel_index2 >= 2097) && (pixel_index2 <= 2103)) || pixel_index2 == 2169 || pixel_index2 == 2177 || ((pixel_index2 >= 2193) && (pixel_index2 <= 2194)) || ((pixel_index2 >= 2198) && (pixel_index2 <= 2199)) || pixel_index2 == 2239 || ((pixel_index2 >= 2241) && (pixel_index2 <= 2242)) || pixel_index2 == 2244 || pixel_index2 == 2247 || pixel_index2 == 2249 || pixel_index2 == 2265 || pixel_index2 == 2273 || ((pixel_index2 >= 2289) && (pixel_index2 <= 2290)) || ((pixel_index2 >= 2294) && (pixel_index2 <= 2295)) || pixel_index2 == 2335 || pixel_index2 == 2337 || pixel_index2 == 2339 || ((pixel_index2 >= 2356) && (pixel_index2 <= 2361)) || ((pixel_index2 >= 2369) && (pixel_index2 <= 2373)) || ((pixel_index2 >= 2385) && (pixel_index2 <= 2391)) || ((pixel_index2 >= 2438) && (pixel_index2 <= 2442)) || ((pixel_index2 >= 2452) && (pixel_index2 <= 2457)) || ((pixel_index2 >= 2465) && (pixel_index2 <= 2469)) || ((pixel_index2 >= 2481) && (pixel_index2 <= 2486)) || pixel_index2 == 2533 || pixel_index2 == 2539 || pixel_index2 == 2549 || ((pixel_index2 >= 2552) && (pixel_index2 <= 2553)) || pixel_index2 == 2561 || ((pixel_index2 >= 2564) && (pixel_index2 <= 2565)) || ((pixel_index2 >= 2627) && (pixel_index2 <= 2629)) || pixel_index2 == 2635 || ((pixel_index2 >= 2637) && (pixel_index2 <= 2638)) || pixel_index2 == 2649 || pixel_index2 == 2657 || ((pixel_index2 >= 2722) && (pixel_index2 <= 2725)) || pixel_index2 == 2731 || ((pixel_index2 >= 2733) && (pixel_index2 <= 2734)) || ((pixel_index2 >= 2743) && (pixel_index2 <= 2755)) || ((pixel_index2 >= 2818) && (pixel_index2 <= 2821)) || pixel_index2 == 2827 || ((pixel_index2 >= 2829) && (pixel_index2 <= 2830)) || ((pixel_index2 >= 2839) && (pixel_index2 <= 2841)) || ((pixel_index2 >= 2849) && (pixel_index2 <= 2851)) || ((pixel_index2 >= 2914) && (pixel_index2 <= 2917)) || pixel_index2 == 2923 || pixel_index2 == 2936 || pixel_index2 == 2945 || pixel_index2 == 2963 || ((pixel_index2 >= 3014) && (pixel_index2 <= 3018)) || ((pixel_index2 >= 3061) && (pixel_index2 <= 3062)) || pixel_index2 == 3064 || ((pixel_index2 >= 3108) && (pixel_index2 <= 3116)) || pixel_index2 == 3160 || ((pixel_index2 >= 3204) && (pixel_index2 <= 3212)) || ((pixel_index2 >= 3300) && (pixel_index2 <= 3308)) || pixel_index2 == 3317 || ((pixel_index2 >= 3319) && (pixel_index2 <= 3320)) || ((pixel_index2 >= 3330) && (pixel_index2 <= 3331)) || pixel_index2 == 3333 || pixel_index2 == 3338 || ((pixel_index2 >= 3396) && (pixel_index2 <= 3404)) || pixel_index2 == 3433 || ((pixel_index2 >= 3436) && (pixel_index2 <= 3437)) || ((pixel_index2 >= 3492) && (pixel_index2 <= 3500)) || ((pixel_index2 >= 3588) && (pixel_index2 <= 3596)) || ((pixel_index2 >= 3684) && (pixel_index2 <= 3692)) || ((pixel_index2 >= 3724) && (pixel_index2 <= 3729)) || ((pixel_index2 >= 3820) && (pixel_index2 <= 3825)) || ((pixel_index2 >= 3893) && (pixel_index2 <= 3894)) || ((pixel_index2 >= 3897) && (pixel_index2 <= 3905)) || ((pixel_index2 >= 3908) && (pixel_index2 <= 3909)) || ((pixel_index2 >= 3989) && (pixel_index2 <= 3990)) || ((pixel_index2 >= 3994) && (pixel_index2 <= 4000)) || ((pixel_index2 >= 4004) && (pixel_index2 <= 4005)) || ((pixel_index2 >= 4085) && (pixel_index2 <= 4086)) || ((pixel_index2 >= 4090) && (pixel_index2 <= 4096)) || ((pixel_index2 >= 4100) && (pixel_index2 <= 4101)) || pixel_index2 == 4706 || pixel_index2 == 4797 || pixel_index2 == 5666 || pixel_index2 == 5757) oled_data2 = 16'b0101001010001010;
                    else if (pixel_index2 == 1296 || ((pixel_index2 >= 1300) && (pixel_index2 <= 1301)) || pixel_index2 == 1303 || pixel_index2 == 1306 || pixel_index2 == 1308 || pixel_index2 == 1310 || pixel_index2 == 1312 || pixel_index2 == 1391 || pixel_index2 == 1396 || pixel_index2 == 1400 || pixel_index2 == 1402 || pixel_index2 == 1405 || ((pixel_index2 >= 1407) && (pixel_index2 <= 1408)) || pixel_index2 == 1489 || ((pixel_index2 >= 1491) && (pixel_index2 <= 1492)) || pixel_index2 == 1494 || pixel_index2 == 1496 || pixel_index2 == 1498 || pixel_index2 == 1501 || pixel_index2 == 1504 || pixel_index2 == 3353 || pixel_index2 == 3449 || pixel_index2 == 3545) oled_data2 = 16'b0101001010010100;
                    else if (((pixel_index2 >= 1317) && (pixel_index2 <= 1319)) || ((pixel_index2 >= 1322) && (pixel_index2 <= 1324)) || ((pixel_index2 >= 1327) && (pixel_index2 <= 1329)) || ((pixel_index2 >= 1332) && (pixel_index2 <= 1334)) || pixel_index2 == 1415 || pixel_index2 == 1420 || pixel_index2 == 1423 || pixel_index2 == 1425 || pixel_index2 == 1430 || ((pixel_index2 >= 1509) && (pixel_index2 <= 1511)) || pixel_index2 == 1516 || pixel_index2 == 1519 || pixel_index2 == 1521 || pixel_index2 == 1526 || pixel_index2 == 1605 || pixel_index2 == 1607 || pixel_index2 == 1612 || pixel_index2 == 1615 || pixel_index2 == 1617 || pixel_index2 == 1622 || pixel_index2 == 1701 || pixel_index2 == 1703 || ((pixel_index2 >= 1706) && (pixel_index2 <= 1708)) || ((pixel_index2 >= 1711) && (pixel_index2 <= 1713)) || (pixel_index2 >= 1716) && (pixel_index2 <= 1718)) oled_data2 = 16'b1010000000001010;
                    else if (((pixel_index2 >= 1578) && (pixel_index2 <= 1582)) || pixel_index2 == 1674 || pixel_index2 == 1678 || pixel_index2 == 1770 || pixel_index2 == 1774 || pixel_index2 == 1866 || pixel_index2 == 1870 || ((pixel_index2 >= 1962) && (pixel_index2 <= 1966)) || pixel_index2 == 2788 || pixel_index2 == 2791 || ((pixel_index2 >= 2794) && (pixel_index2 <= 2795)) || ((pixel_index2 >= 2799) && (pixel_index2 <= 2800)) || ((pixel_index2 >= 2804) && (pixel_index2 <= 2805)) || pixel_index2 == 2885 || pixel_index2 == 2887 || pixel_index2 == 2889 || pixel_index2 == 2892 || pixel_index2 == 2894 || pixel_index2 == 2897 || pixel_index2 == 2899 || pixel_index2 == 2902 || pixel_index2 == 2905 || ((pixel_index2 >= 2982) && (pixel_index2 <= 2983)) || pixel_index2 == 2988 || pixel_index2 == 2990 || pixel_index2 == 2993 || pixel_index2 == 2998 || pixel_index2 == 3000 || pixel_index2 == 3077 || pixel_index2 == 3079 || pixel_index2 == 3081 || pixel_index2 == 3084 || pixel_index2 == 3086 || pixel_index2 == 3089 || pixel_index2 == 3091 || pixel_index2 == 3094 || pixel_index2 == 3097 || pixel_index2 == 3172 || pixel_index2 == 3175 || ((pixel_index2 >= 3178) && (pixel_index2 <= 3179)) || ((pixel_index2 >= 3183) && (pixel_index2 <= 3184)) || (pixel_index2 >= 3188) && (pixel_index2 <= 3189)) oled_data2 = 16'b1111010100001010;
                    else if (pixel_index2 == 3229 || (pixel_index2 >= 3325) && (pixel_index2 <= 3326)) oled_data2 = 16'b0101010100001010;
                    else if (pixel_index2 == 3394 || pixel_index2 == 3490) oled_data2 = 16'b0000000000010100;
                    else if (pixel_index2 == 3532 || pixel_index2 == 3537) oled_data2 = 16'b0101000000000000;
                    else if (((pixel_index2 >= 4423) && (pixel_index2 <= 4505)) || ((pixel_index2 >= 4513) && (pixel_index2 <= 4518)) || (pixel_index2 >= 4602) && (pixel_index2 <= 4606)) oled_data2 = 16'b0000001010011110;
                    else if (((pixel_index2 >= 4519) && (pixel_index2 <= 4601)) || ((pixel_index2 >= 4609) && (pixel_index2 <= 4619)) || ((pixel_index2 >= 4693) && (pixel_index2 <= 4702)) || pixel_index2 == 4705 || pixel_index2 == 4798 || pixel_index2 == 4801 || pixel_index2 == 4894 || ((pixel_index2 >= 4897) && (pixel_index2 <= 4898)) || ((pixel_index2 >= 4989) && (pixel_index2 <= 4990)) || pixel_index2 == 4993 || pixel_index2 == 5086 || pixel_index2 == 5089 || pixel_index2 == 5182 || pixel_index2 == 5185 || pixel_index2 == 5278 || pixel_index2 == 5281 || pixel_index2 == 5374 || pixel_index2 == 5377 || pixel_index2 == 5470 || pixel_index2 == 5473 || pixel_index2 == 5566 || pixel_index2 == 5569 || pixel_index2 == 5662 || pixel_index2 == 5665 || pixel_index2 == 5758 || pixel_index2 == 5761 || pixel_index2 == 5854 || ((pixel_index2 >= 5857) && (pixel_index2 <= 5867)) || ((pixel_index2 >= 5941) && (pixel_index2 <= 5950)) || (pixel_index2 >= 5959) && (pixel_index2 <= 6041)) oled_data2 = 16'b0000001010010100;
                    else if (pixel_index2 == 4813 || pixel_index2 == 4818 || ((pixel_index2 >= 4821) && (pixel_index2 <= 4826)) || ((pixel_index2 >= 4830) && (pixel_index2 <= 4833)) || ((pixel_index2 >= 4836) && (pixel_index2 <= 4837)) || pixel_index2 == 4840 || pixel_index2 == 4844 || ((pixel_index2 >= 4847) && (pixel_index2 <= 4850)) || pixel_index2 == 4862 || ((pixel_index2 >= 4866) && (pixel_index2 <= 4867)) || pixel_index2 == 4870 || ((pixel_index2 >= 4874) && (pixel_index2 <= 4879)) || ((pixel_index2 >= 4883) && (pixel_index2 <= 4886)) || pixel_index2 == 4908 || pixel_index2 == 4913 || pixel_index2 == 4916 || pixel_index2 == 4923 || pixel_index2 == 4925 || pixel_index2 == 4930 || pixel_index2 == 4934 || pixel_index2 == 4937 || pixel_index2 == 4939 || pixel_index2 == 4942 || pixel_index2 == 4947 || pixel_index2 == 4957 || pixel_index2 == 4964 || pixel_index2 == 4967 || pixel_index2 == 4969 || pixel_index2 == 4976 || pixel_index2 == 4978 || pixel_index2 == 4983 || pixel_index2 == 5031 || pixel_index2 == 5061 || pixel_index2 == 5221 || pixel_index2 == 5251 || ((pixel_index2 >= 5268) && (pixel_index2 <= 5270)) || pixel_index2 == 5316 || pixel_index2 == 5346 || pixel_index2 == 5367 || pixel_index2 == 5504 || pixel_index2 == 5521 || pixel_index2 == 5547 || pixel_index2 == 5550 || pixel_index2 == 5557 || ((pixel_index2 >= 5576) && (pixel_index2 <= 5579)) || ((pixel_index2 >= 5582) && (pixel_index2 <= 5583)) || ((pixel_index2 >= 5597) && (pixel_index2 <= 5599)) || ((pixel_index2 >= 5606) && (pixel_index2 <= 5607)) || ((pixel_index2 >= 5614) && (pixel_index2 <= 5616)) || ((pixel_index2 >= 5625) && (pixel_index2 <= 5628)) || ((pixel_index2 >= 5631) && (pixel_index2 <= 5632)) || ((pixel_index2 >= 5636) && (pixel_index2 <= 5637)) || ((pixel_index2 >= 5644) && (pixel_index2 <= 5645)) || (pixel_index2 >= 5650) && (pixel_index2 <= 5652)) oled_data2 = 16'b0101001010000000;
                    else if (pixel_index2 == 4909 || pixel_index2 == 4914 || ((pixel_index2 >= 4917) && (pixel_index2 <= 4922)) || ((pixel_index2 >= 4926) && (pixel_index2 <= 4929)) || ((pixel_index2 >= 4932) && (pixel_index2 <= 4933)) || pixel_index2 == 4936 || pixel_index2 == 4940 || ((pixel_index2 >= 4943) && (pixel_index2 <= 4946)) || pixel_index2 == 4958 || ((pixel_index2 >= 4962) && (pixel_index2 <= 4963)) || pixel_index2 == 4966 || ((pixel_index2 >= 4970) && (pixel_index2 <= 4975)) || ((pixel_index2 >= 4979) && (pixel_index2 <= 4982)) || ((pixel_index2 >= 5004) && (pixel_index2 <= 5005)) || ((pixel_index2 >= 5009) && (pixel_index2 <= 5010)) || ((pixel_index2 >= 5012) && (pixel_index2 <= 5019)) || ((pixel_index2 >= 5021) && (pixel_index2 <= 5026)) || ((pixel_index2 >= 5028) && (pixel_index2 <= 5030)) || ((pixel_index2 >= 5032) && (pixel_index2 <= 5033)) || ((pixel_index2 >= 5035) && (pixel_index2 <= 5036)) || ((pixel_index2 >= 5038) && (pixel_index2 <= 5043)) || ((pixel_index2 >= 5053) && (pixel_index2 <= 5054)) || ((pixel_index2 >= 5058) && (pixel_index2 <= 5060)) || ((pixel_index2 >= 5062) && (pixel_index2 <= 5063)) || ((pixel_index2 >= 5065) && (pixel_index2 <= 5072)) || ((pixel_index2 >= 5074) && (pixel_index2 <= 5079)) || ((pixel_index2 >= 5100) && (pixel_index2 <= 5101)) || ((pixel_index2 >= 5105) && (pixel_index2 <= 5106)) || ((pixel_index2 >= 5108) && (pixel_index2 <= 5110)) || ((pixel_index2 >= 5113) && (pixel_index2 <= 5115)) || ((pixel_index2 >= 5120) && (pixel_index2 <= 5122)) || ((pixel_index2 >= 5125) && (pixel_index2 <= 5129)) || ((pixel_index2 >= 5131) && (pixel_index2 <= 5132)) || ((pixel_index2 >= 5137) && (pixel_index2 <= 5139)) || ((pixel_index2 >= 5149) && (pixel_index2 <= 5150)) || ((pixel_index2 >= 5155) && (pixel_index2 <= 5159)) || ((pixel_index2 >= 5161) && (pixel_index2 <= 5163)) || ((pixel_index2 >= 5166) && (pixel_index2 <= 5168)) || ((pixel_index2 >= 5170) && (pixel_index2 <= 5172)) || ((pixel_index2 >= 5196) && (pixel_index2 <= 5197)) || ((pixel_index2 >= 5201) && (pixel_index2 <= 5202)) || ((pixel_index2 >= 5204) && (pixel_index2 <= 5205)) || ((pixel_index2 >= 5210) && (pixel_index2 <= 5211)) || ((pixel_index2 >= 5217) && (pixel_index2 <= 5218)) || ((pixel_index2 >= 5222) && (pixel_index2 <= 5225)) || ((pixel_index2 >= 5227) && (pixel_index2 <= 5228)) || ((pixel_index2 >= 5234) && (pixel_index2 <= 5235)) || ((pixel_index2 >= 5245) && (pixel_index2 <= 5246)) || ((pixel_index2 >= 5252) && (pixel_index2 <= 5255)) || ((pixel_index2 >= 5257) && (pixel_index2 <= 5258)) || ((pixel_index2 >= 5263) && (pixel_index2 <= 5264)) || ((pixel_index2 >= 5266) && (pixel_index2 <= 5267)) || ((pixel_index2 >= 5292) && (pixel_index2 <= 5293)) || ((pixel_index2 >= 5297) && (pixel_index2 <= 5298)) || ((pixel_index2 >= 5300) && (pixel_index2 <= 5301)) || ((pixel_index2 >= 5306) && (pixel_index2 <= 5307)) || ((pixel_index2 >= 5313) && (pixel_index2 <= 5314)) || ((pixel_index2 >= 5317) && (pixel_index2 <= 5321)) || ((pixel_index2 >= 5323) && (pixel_index2 <= 5324)) || ((pixel_index2 >= 5330) && (pixel_index2 <= 5331)) || ((pixel_index2 >= 5341) && (pixel_index2 <= 5342)) || ((pixel_index2 >= 5347) && (pixel_index2 <= 5351)) || ((pixel_index2 >= 5353) && (pixel_index2 <= 5354)) || ((pixel_index2 >= 5359) && (pixel_index2 <= 5360)) || ((pixel_index2 >= 5362) && (pixel_index2 <= 5366)) || ((pixel_index2 >= 5388) && (pixel_index2 <= 5389)) || ((pixel_index2 >= 5393) && (pixel_index2 <= 5394)) || ((pixel_index2 >= 5396) && (pixel_index2 <= 5397)) || ((pixel_index2 >= 5402) && (pixel_index2 <= 5403)) || ((pixel_index2 >= 5409) && (pixel_index2 <= 5410)) || ((pixel_index2 >= 5412) && (pixel_index2 <= 5414)) || ((pixel_index2 >= 5416) && (pixel_index2 <= 5417)) || ((pixel_index2 >= 5419) && (pixel_index2 <= 5420)) || ((pixel_index2 >= 5426) && (pixel_index2 <= 5427)) || ((pixel_index2 >= 5437) && (pixel_index2 <= 5438)) || ((pixel_index2 >= 5442) && (pixel_index2 <= 5444)) || ((pixel_index2 >= 5446) && (pixel_index2 <= 5447)) || ((pixel_index2 >= 5449) && (pixel_index2 <= 5450)) || ((pixel_index2 >= 5455) && (pixel_index2 <= 5456)) || ((pixel_index2 >= 5459) && (pixel_index2 <= 5463)) || ((pixel_index2 >= 5484) && (pixel_index2 <= 5485)) || ((pixel_index2 >= 5489) && (pixel_index2 <= 5490)) || ((pixel_index2 >= 5492) && (pixel_index2 <= 5493)) || ((pixel_index2 >= 5498) && (pixel_index2 <= 5499)) || ((pixel_index2 >= 5505) && (pixel_index2 <= 5506)) || ((pixel_index2 >= 5508) && (pixel_index2 <= 5509)) || ((pixel_index2 >= 5512) && (pixel_index2 <= 5513)) || ((pixel_index2 >= 5515) && (pixel_index2 <= 5516)) || ((pixel_index2 >= 5522) && (pixel_index2 <= 5523)) || ((pixel_index2 >= 5533) && (pixel_index2 <= 5534)) || ((pixel_index2 >= 5538) && (pixel_index2 <= 5539)) || ((pixel_index2 >= 5542) && (pixel_index2 <= 5543)) || ((pixel_index2 >= 5545) && (pixel_index2 <= 5546)) || ((pixel_index2 >= 5551) && (pixel_index2 <= 5552)) || ((pixel_index2 >= 5558) && (pixel_index2 <= 5559)) || ((pixel_index2 >= 5580) && (pixel_index2 <= 5581)) || ((pixel_index2 >= 5585) && (pixel_index2 <= 5586)) || ((pixel_index2 >= 5588) && (pixel_index2 <= 5589)) || ((pixel_index2 >= 5594) && (pixel_index2 <= 5595)) || ((pixel_index2 >= 5600) && (pixel_index2 <= 5602)) || ((pixel_index2 >= 5604) && (pixel_index2 <= 5605)) || ((pixel_index2 >= 5608) && (pixel_index2 <= 5609)) || ((pixel_index2 >= 5611) && (pixel_index2 <= 5612)) || ((pixel_index2 >= 5617) && (pixel_index2 <= 5619)) || ((pixel_index2 >= 5629) && (pixel_index2 <= 5630)) || ((pixel_index2 >= 5634) && (pixel_index2 <= 5635)) || ((pixel_index2 >= 5638) && (pixel_index2 <= 5639)) || ((pixel_index2 >= 5641) && (pixel_index2 <= 5643)) || ((pixel_index2 >= 5646) && (pixel_index2 <= 5648)) || ((pixel_index2 >= 5653) && (pixel_index2 <= 5655)) || ((pixel_index2 >= 5672) && (pixel_index2 <= 5679)) || ((pixel_index2 >= 5681) && (pixel_index2 <= 5682)) || ((pixel_index2 >= 5684) && (pixel_index2 <= 5685)) || ((pixel_index2 >= 5690) && (pixel_index2 <= 5691)) || ((pixel_index2 >= 5693) && (pixel_index2 <= 5698)) || ((pixel_index2 >= 5700) && (pixel_index2 <= 5705)) || ((pixel_index2 >= 5707) && (pixel_index2 <= 5708)) || ((pixel_index2 >= 5710) && (pixel_index2 <= 5715)) || ((pixel_index2 >= 5721) && (pixel_index2 <= 5728)) || ((pixel_index2 >= 5730) && (pixel_index2 <= 5735)) || ((pixel_index2 >= 5737) && (pixel_index2 <= 5744)) || ((pixel_index2 >= 5746) && (pixel_index2 <= 5751)) || ((pixel_index2 >= 5769) && (pixel_index2 <= 5774)) || pixel_index2 == 5777 || pixel_index2 == 5781 || pixel_index2 == 5786 || ((pixel_index2 >= 5790) && (pixel_index2 <= 5793)) || ((pixel_index2 >= 5797) && (pixel_index2 <= 5800)) || pixel_index2 == 5803 || ((pixel_index2 >= 5807) && (pixel_index2 <= 5810)) || ((pixel_index2 >= 5818) && (pixel_index2 <= 5823)) || ((pixel_index2 >= 5827) && (pixel_index2 <= 5830)) || ((pixel_index2 >= 5834) && (pixel_index2 <= 5839)) || (pixel_index2 >= 5843) && (pixel_index2 <= 5846)) oled_data2 = 16'b1111010100010100;
                    else oled_data2 = 0;
                end
                5: begin
                    if (pixel_index2 == 97 || pixel_index2 == 99 || pixel_index2 == 101 || ((pixel_index2 >= 103) && (pixel_index2 <= 104)) || ((pixel_index2 >= 106) && (pixel_index2 <= 109)) || pixel_index2 == 111 || ((pixel_index2 >= 113) && (pixel_index2 <= 114)) || ((pixel_index2 >= 118) && (pixel_index2 <= 120)) || pixel_index2 == 195 || pixel_index2 == 197 || ((pixel_index2 >= 199) && (pixel_index2 <= 200)) || pixel_index2 == 202 || ((pixel_index2 >= 204) && (pixel_index2 <= 205)) || pixel_index2 == 207 || ((pixel_index2 >= 209) && (pixel_index2 <= 210)) || pixel_index2 == 213 || pixel_index2 == 289 || ((pixel_index2 >= 291) && (pixel_index2 <= 296)) || pixel_index2 == 298 || ((pixel_index2 >= 300) && (pixel_index2 <= 301)) || pixel_index2 == 303 || ((pixel_index2 >= 305) && (pixel_index2 <= 306)) || ((pixel_index2 >= 310) && (pixel_index2 <= 312)) || pixel_index2 == 385 || ((pixel_index2 >= 387) && (pixel_index2 <= 392)) || pixel_index2 == 394 || ((pixel_index2 >= 396) && (pixel_index2 <= 397)) || ((pixel_index2 >= 399) && (pixel_index2 <= 402)) || pixel_index2 == 408 || ((pixel_index2 >= 501) && (pixel_index2 <= 504)) || ((pixel_index2 >= 674) && (pixel_index2 <= 675)) || ((pixel_index2 >= 678) && (pixel_index2 <= 681)) || ((pixel_index2 >= 685) && (pixel_index2 <= 686)) || pixel_index2 == 688 || ((pixel_index2 >= 690) && (pixel_index2 <= 691)) || ((pixel_index2 >= 693) && (pixel_index2 <= 696)) || ((pixel_index2 >= 770) && (pixel_index2 <= 771)) || pixel_index2 == 774 || ((pixel_index2 >= 776) && (pixel_index2 <= 777)) || ((pixel_index2 >= 779) && (pixel_index2 <= 782)) || pixel_index2 == 784 || ((pixel_index2 >= 786) && (pixel_index2 <= 787)) || ((pixel_index2 >= 790) && (pixel_index2 <= 791)) || ((pixel_index2 >= 866) && (pixel_index2 <= 867)) || pixel_index2 == 870 || ((pixel_index2 >= 872) && (pixel_index2 <= 873)) || pixel_index2 == 875 || ((pixel_index2 >= 877) && (pixel_index2 <= 878)) || pixel_index2 == 880 || ((pixel_index2 >= 882) && (pixel_index2 <= 883)) || ((pixel_index2 >= 886) && (pixel_index2 <= 887)) || ((pixel_index2 >= 895) && (pixel_index2 <= 896)) || ((pixel_index2 >= 899) && (pixel_index2 <= 900)) || ((pixel_index2 >= 903) && (pixel_index2 <= 904)) || ((pixel_index2 >= 907) && (pixel_index2 <= 908)) || ((pixel_index2 >= 911) && (pixel_index2 <= 912)) || ((pixel_index2 >= 915) && (pixel_index2 <= 916)) || ((pixel_index2 >= 919) && (pixel_index2 <= 920)) || ((pixel_index2 >= 923) && (pixel_index2 <= 924)) || ((pixel_index2 >= 927) && (pixel_index2 <= 928)) || ((pixel_index2 >= 931) && (pixel_index2 <= 932)) || ((pixel_index2 >= 935) && (pixel_index2 <= 936)) || ((pixel_index2 >= 939) && (pixel_index2 <= 940)) || ((pixel_index2 >= 943) && (pixel_index2 <= 944)) || ((pixel_index2 >= 947) && (pixel_index2 <= 948)) || ((pixel_index2 >= 951) && (pixel_index2 <= 952)) || ((pixel_index2 >= 955) && (pixel_index2 <= 956)) || ((pixel_index2 >= 961) && (pixel_index2 <= 964)) || pixel_index2 == 966 || ((pixel_index2 >= 968) && (pixel_index2 <= 969)) || ((pixel_index2 >= 971) && (pixel_index2 <= 974)) || ((pixel_index2 >= 976) && (pixel_index2 <= 979)) || ((pixel_index2 >= 981) && (pixel_index2 <= 984)) || ((pixel_index2 >= 1637) && (pixel_index2 <= 1638)) || ((pixel_index2 >= 1641) && (pixel_index2 <= 1644)) || ((pixel_index2 >= 1646) && (pixel_index2 <= 1649)) || ((pixel_index2 >= 1652) && (pixel_index2 <= 1654)) || pixel_index2 == 1732 || pixel_index2 == 1735 || pixel_index2 == 1740 || pixel_index2 == 1745 || pixel_index2 == 1747 || pixel_index2 == 1831 || pixel_index2 == 1836 || ((pixel_index2 >= 1839) && (pixel_index2 <= 1841)) || ((pixel_index2 >= 1844) && (pixel_index2 <= 1845)) || pixel_index2 == 1924 || pixel_index2 == 1927 || pixel_index2 == 1932 || pixel_index2 == 1937 || pixel_index2 == 1942 || ((pixel_index2 >= 2021) && (pixel_index2 <= 2022)) || pixel_index2 == 2028 || ((pixel_index2 >= 2030) && (pixel_index2 <= 2033)) || ((pixel_index2 >= 2035) && (pixel_index2 <= 2037)) || pixel_index2 == 2788 || pixel_index2 == 2791 || ((pixel_index2 >= 2794) && (pixel_index2 <= 2795)) || ((pixel_index2 >= 2799) && (pixel_index2 <= 2800)) || ((pixel_index2 >= 2804) && (pixel_index2 <= 2805)) || pixel_index2 == 2885 || pixel_index2 == 2887 || pixel_index2 == 2889 || pixel_index2 == 2892 || pixel_index2 == 2894 || pixel_index2 == 2897 || pixel_index2 == 2899 || pixel_index2 == 2902 || ((pixel_index2 >= 2982) && (pixel_index2 <= 2983)) || pixel_index2 == 2988 || pixel_index2 == 2990 || pixel_index2 == 2993 || pixel_index2 == 2998 || pixel_index2 == 3077 || pixel_index2 == 3079 || pixel_index2 == 3081 || pixel_index2 == 3084 || pixel_index2 == 3086 || pixel_index2 == 3089 || pixel_index2 == 3091 || pixel_index2 == 3094 || ((pixel_index2 >= 3133) && (pixel_index2 <= 3134)) || pixel_index2 == 3172 || pixel_index2 == 3175 || ((pixel_index2 >= 3178) && (pixel_index2 <= 3179)) || ((pixel_index2 >= 3183) && (pixel_index2 <= 3184)) || ((pixel_index2 >= 3188) && (pixel_index2 <= 3189)) || pixel_index2 == 3228 || pixel_index2 == 3327 || ((pixel_index2 >= 3364) && (pixel_index2 <= 3367)) || ((pixel_index2 >= 3370) && (pixel_index2 <= 3372)) || ((pixel_index2 >= 3375) && (pixel_index2 <= 3376)) || ((pixel_index2 >= 3380) && (pixel_index2 <= 3382)) || pixel_index2 == 3463 || pixel_index2 == 3465 || pixel_index2 == 3468 || pixel_index2 == 3470 || pixel_index2 == 3473 || pixel_index2 == 3475 || pixel_index2 == 3478 || pixel_index2 == 3559 || ((pixel_index2 >= 3562) && (pixel_index2 <= 3564)) || pixel_index2 == 3566 || pixel_index2 == 3569 || ((pixel_index2 >= 3572) && (pixel_index2 <= 3574)) || ((pixel_index2 >= 3630) && (pixel_index2 <= 3631)) || pixel_index2 == 3655 || pixel_index2 == 3657 || pixel_index2 == 3660 || pixel_index2 == 3662 || pixel_index2 == 3665 || pixel_index2 == 3667 || pixel_index2 == 3670 || pixel_index2 == 3751 || ((pixel_index2 >= 3754) && (pixel_index2 <= 3756)) || pixel_index2 == 3758 || pixel_index2 == 3761 || ((pixel_index2 >= 3764) && (pixel_index2 <= 3766)) || ((pixel_index2 >= 3938) && (pixel_index2 <= 3939)) || pixel_index2 == 3942 || pixel_index2 == 3945 || ((pixel_index2 >= 3947) && (pixel_index2 <= 3950)) || pixel_index2 == 3952 || ((pixel_index2 >= 3954) && (pixel_index2 <= 3955)) || ((pixel_index2 >= 3959) && (pixel_index2 <= 3962)) || ((pixel_index2 >= 3964) && (pixel_index2 <= 3967)) || ((pixel_index2 >= 3969) && (pixel_index2 <= 3972)) || ((pixel_index2 >= 3974) && (pixel_index2 <= 3977)) || pixel_index2 == 3979 || ((pixel_index2 >= 3981) && (pixel_index2 <= 3982)) || ((pixel_index2 >= 3984) && (pixel_index2 <= 3986)) || ((pixel_index2 >= 4034) && (pixel_index2 <= 4035)) || ((pixel_index2 >= 4039) && (pixel_index2 <= 4040)) || ((pixel_index2 >= 4045) && (pixel_index2 <= 4046)) || pixel_index2 == 4048 || ((pixel_index2 >= 4050) && (pixel_index2 <= 4051)) || ((pixel_index2 >= 4057) && (pixel_index2 <= 4058)) || ((pixel_index2 >= 4060) && (pixel_index2 <= 4061)) || pixel_index2 == 4065 || ((pixel_index2 >= 4067) && (pixel_index2 <= 4068)) || pixel_index2 == 4070 || ((pixel_index2 >= 4072) && (pixel_index2 <= 4073)) || ((pixel_index2 >= 4075) && (pixel_index2 <= 4078)) || ((pixel_index2 >= 4082) && (pixel_index2 <= 4083)) || ((pixel_index2 >= 4130) && (pixel_index2 <= 4131)) || ((pixel_index2 >= 4135) && (pixel_index2 <= 4136)) || ((pixel_index2 >= 4139) && (pixel_index2 <= 4140)) || pixel_index2 == 4142 || pixel_index2 == 4144 || ((pixel_index2 >= 4146) && (pixel_index2 <= 4147)) || ((pixel_index2 >= 4151) && (pixel_index2 <= 4152)) || pixel_index2 == 4154 || ((pixel_index2 >= 4157) && (pixel_index2 <= 4159)) || pixel_index2 == 4161 || ((pixel_index2 >= 4163) && (pixel_index2 <= 4164)) || pixel_index2 == 4166 || ((pixel_index2 >= 4168) && (pixel_index2 <= 4169)) || pixel_index2 == 4171 || ((pixel_index2 >= 4173) && (pixel_index2 <= 4174)) || ((pixel_index2 >= 4178) && (pixel_index2 <= 4179)) || ((pixel_index2 >= 4225) && (pixel_index2 <= 4228)) || pixel_index2 == 4230 || pixel_index2 == 4233 || ((pixel_index2 >= 4235) && (pixel_index2 <= 4238)) || ((pixel_index2 >= 4240) && (pixel_index2 <= 4243)) || ((pixel_index2 >= 4247) && (pixel_index2 <= 4250)) || ((pixel_index2 >= 4252) && (pixel_index2 <= 4254)) || ((pixel_index2 >= 4257) && (pixel_index2 <= 4260)) || ((pixel_index2 >= 4262) && (pixel_index2 <= 4265)) || pixel_index2 == 4267 || ((pixel_index2 >= 4269) && (pixel_index2 <= 4270)) || ((pixel_index2 >= 4272) && (pixel_index2 <= 4274)) || pixel_index2 == 4802 || pixel_index2 == 4893 || pixel_index2 == 5762 || pixel_index2 == 5853) oled_data2 = 16'b1111011110011110;
                    else if (pixel_index2 == 124 || ((pixel_index2 >= 130) && (pixel_index2 <= 184)) || pixel_index2 == 190 || pixel_index2 == 220 || pixel_index2 == 229 || pixel_index2 == 233 || pixel_index2 == 237 || pixel_index2 == 241 || pixel_index2 == 245 || pixel_index2 == 249 || pixel_index2 == 253 || pixel_index2 == 257 || pixel_index2 == 261 || pixel_index2 == 265 || pixel_index2 == 269 || pixel_index2 == 273 || pixel_index2 == 277 || pixel_index2 == 286 || pixel_index2 == 316 || pixel_index2 == 325 || pixel_index2 == 329 || pixel_index2 == 333 || pixel_index2 == 337 || pixel_index2 == 341 || pixel_index2 == 345 || pixel_index2 == 349 || pixel_index2 == 353 || pixel_index2 == 357 || pixel_index2 == 361 || pixel_index2 == 365 || pixel_index2 == 369 || pixel_index2 == 373 || pixel_index2 == 382 || pixel_index2 == 412 || pixel_index2 == 421 || pixel_index2 == 425 || pixel_index2 == 429 || pixel_index2 == 433 || pixel_index2 == 437 || pixel_index2 == 441 || pixel_index2 == 445 || pixel_index2 == 449 || pixel_index2 == 453 || pixel_index2 == 457 || pixel_index2 == 461 || pixel_index2 == 465 || pixel_index2 == 469 || pixel_index2 == 478 || pixel_index2 == 508 || pixel_index2 == 517 || pixel_index2 == 521 || pixel_index2 == 525 || pixel_index2 == 529 || pixel_index2 == 533 || pixel_index2 == 537 || pixel_index2 == 541 || pixel_index2 == 545 || pixel_index2 == 549 || pixel_index2 == 553 || pixel_index2 == 557 || pixel_index2 == 561 || pixel_index2 == 565 || pixel_index2 == 574 || pixel_index2 == 604 || pixel_index2 == 613 || pixel_index2 == 617 || pixel_index2 == 621 || pixel_index2 == 625 || pixel_index2 == 629 || pixel_index2 == 633 || pixel_index2 == 637 || pixel_index2 == 641 || pixel_index2 == 645 || pixel_index2 == 649 || pixel_index2 == 653 || pixel_index2 == 657 || pixel_index2 == 661 || pixel_index2 == 670 || pixel_index2 == 700 || pixel_index2 == 709 || pixel_index2 == 713 || pixel_index2 == 717 || pixel_index2 == 721 || pixel_index2 == 725 || pixel_index2 == 729 || pixel_index2 == 733 || pixel_index2 == 737 || pixel_index2 == 741 || pixel_index2 == 745 || pixel_index2 == 749 || pixel_index2 == 753 || pixel_index2 == 757 || pixel_index2 == 766 || pixel_index2 == 796 || ((pixel_index2 >= 802) && (pixel_index2 <= 856)) || pixel_index2 == 862 || ((pixel_index2 >= 892) && (pixel_index2 <= 894)) || ((pixel_index2 >= 897) && (pixel_index2 <= 898)) || ((pixel_index2 >= 901) && (pixel_index2 <= 902)) || ((pixel_index2 >= 905) && (pixel_index2 <= 906)) || ((pixel_index2 >= 909) && (pixel_index2 <= 910)) || ((pixel_index2 >= 913) && (pixel_index2 <= 914)) || ((pixel_index2 >= 917) && (pixel_index2 <= 918)) || ((pixel_index2 >= 921) && (pixel_index2 <= 922)) || ((pixel_index2 >= 925) && (pixel_index2 <= 926)) || ((pixel_index2 >= 929) && (pixel_index2 <= 930)) || ((pixel_index2 >= 933) && (pixel_index2 <= 934)) || ((pixel_index2 >= 937) && (pixel_index2 <= 938)) || ((pixel_index2 >= 941) && (pixel_index2 <= 942)) || ((pixel_index2 >= 945) && (pixel_index2 <= 946)) || ((pixel_index2 >= 949) && (pixel_index2 <= 950)) || ((pixel_index2 >= 953) && (pixel_index2 <= 954)) || ((pixel_index2 >= 957) && (pixel_index2 <= 958)) || ((pixel_index2 >= 988) && (pixel_index2 <= 1054)) || ((pixel_index2 >= 1084) && (pixel_index2 <= 1085)) || ((pixel_index2 >= 1087) && (pixel_index2 <= 1089)) || ((pixel_index2 >= 1091) && (pixel_index2 <= 1093)) || ((pixel_index2 >= 1095) && (pixel_index2 <= 1097)) || ((pixel_index2 >= 1099) && (pixel_index2 <= 1101)) || ((pixel_index2 >= 1103) && (pixel_index2 <= 1105)) || ((pixel_index2 >= 1107) && (pixel_index2 <= 1109)) || ((pixel_index2 >= 1111) && (pixel_index2 <= 1113)) || ((pixel_index2 >= 1115) && (pixel_index2 <= 1117)) || ((pixel_index2 >= 1119) && (pixel_index2 <= 1121)) || ((pixel_index2 >= 1123) && (pixel_index2 <= 1125)) || ((pixel_index2 >= 1127) && (pixel_index2 <= 1129)) || ((pixel_index2 >= 1131) && (pixel_index2 <= 1133)) || ((pixel_index2 >= 1135) && (pixel_index2 <= 1137)) || ((pixel_index2 >= 1139) && (pixel_index2 <= 1141)) || ((pixel_index2 >= 1143) && (pixel_index2 <= 1145)) || ((pixel_index2 >= 1147) && (pixel_index2 <= 1150)) || ((pixel_index2 >= 1182) && (pixel_index2 <= 1219)) || ((pixel_index2 >= 1240) && (pixel_index2 <= 1244)) || ((pixel_index2 >= 1278) && (pixel_index2 <= 1280)) || ((pixel_index2 >= 1283) && (pixel_index2 <= 1286)) || ((pixel_index2 >= 1290) && (pixel_index2 <= 1291)) || ((pixel_index2 >= 1293) && (pixel_index2 <= 1294)) || ((pixel_index2 >= 1314) && (pixel_index2 <= 1315)) || ((pixel_index2 >= 1336) && (pixel_index2 <= 1340)) || ((pixel_index2 >= 1374) && (pixel_index2 <= 1376)) || ((pixel_index2 >= 1378) && (pixel_index2 <= 1382)) || ((pixel_index2 >= 1386) && (pixel_index2 <= 1390)) || ((pixel_index2 >= 1410) && (pixel_index2 <= 1411)) || ((pixel_index2 >= 1432) && (pixel_index2 <= 1436)) || ((pixel_index2 >= 1470) && (pixel_index2 <= 1478)) || ((pixel_index2 >= 1482) && (pixel_index2 <= 1486)) || ((pixel_index2 >= 1506) && (pixel_index2 <= 1507)) || ((pixel_index2 >= 1528) && (pixel_index2 <= 1532)) || ((pixel_index2 >= 1566) && (pixel_index2 <= 1569)) || ((pixel_index2 >= 1575) && (pixel_index2 <= 1603)) || ((pixel_index2 >= 1624) && (pixel_index2 <= 1628)) || ((pixel_index2 >= 1662) && (pixel_index2 <= 1665)) || pixel_index2 == 1674 || ((pixel_index2 >= 1678) && (pixel_index2 <= 1696)) || ((pixel_index2 >= 1698) && (pixel_index2 <= 1699)) || ((pixel_index2 >= 1720) && (pixel_index2 <= 1724)) || ((pixel_index2 >= 1758) && (pixel_index2 <= 1761)) || pixel_index2 == 1770 || ((pixel_index2 >= 1774) && (pixel_index2 <= 1775)) || ((pixel_index2 >= 1777) && (pixel_index2 <= 1789)) || pixel_index2 == 1792 || ((pixel_index2 >= 1794) && (pixel_index2 <= 1795)) || pixel_index2 == 1816 || ((pixel_index2 >= 1818) && (pixel_index2 <= 1820)) || ((pixel_index2 >= 1854) && (pixel_index2 <= 1857)) || pixel_index2 == 1866 || pixel_index2 == 1870 || ((pixel_index2 >= 1872) && (pixel_index2 <= 1878)) || ((pixel_index2 >= 1882) && (pixel_index2 <= 1888)) || ((pixel_index2 >= 1892) && (pixel_index2 <= 1913)) || ((pixel_index2 >= 1915) && (pixel_index2 <= 1916)) || ((pixel_index2 >= 1948) && (pixel_index2 <= 1953)) || ((pixel_index2 >= 1959) && (pixel_index2 <= 1973)) || pixel_index2 == 1988 || pixel_index2 == 1991 || ((pixel_index2 >= 1993) && (pixel_index2 <= 1994)) || pixel_index2 == 1996 || ((pixel_index2 >= 2000) && (pixel_index2 <= 2001)) || pixel_index2 == 2008 || ((pixel_index2 >= 2011) && (pixel_index2 <= 2014)) || ((pixel_index2 >= 2044) && (pixel_index2 <= 2046)) || ((pixel_index2 >= 2048) && (pixel_index2 <= 2054)) || ((pixel_index2 >= 2058) && (pixel_index2 <= 2069)) || ((pixel_index2 >= 2084) && (pixel_index2 <= 2085)) || pixel_index2 == 2089 || ((pixel_index2 >= 2091) && (pixel_index2 <= 2093)) || ((pixel_index2 >= 2095) && (pixel_index2 <= 2096)) || ((pixel_index2 >= 2104) && (pixel_index2 <= 2105)) || ((pixel_index2 >= 2107) && (pixel_index2 <= 2110)) || pixel_index2 == 2140 || pixel_index2 == 2142 || ((pixel_index2 >= 2144) && (pixel_index2 <= 2150)) || pixel_index2 == 2154 || ((pixel_index2 >= 2157) && (pixel_index2 <= 2168)) || pixel_index2 == 2178 || ((pixel_index2 >= 2180) && (pixel_index2 <= 2184)) || pixel_index2 == 2188 || ((pixel_index2 >= 2190) && (pixel_index2 <= 2192)) || ((pixel_index2 >= 2195) && (pixel_index2 <= 2197)) || ((pixel_index2 >= 2200) && (pixel_index2 <= 2206)) || ((pixel_index2 >= 2236) && (pixel_index2 <= 2238)) || ((pixel_index2 >= 2245) && (pixel_index2 <= 2246)) || pixel_index2 == 2250 || ((pixel_index2 >= 2252) && (pixel_index2 <= 2264)) || ((pixel_index2 >= 2274) && (pixel_index2 <= 2288)) || ((pixel_index2 >= 2291) && (pixel_index2 <= 2293)) || ((pixel_index2 >= 2296) && (pixel_index2 <= 2302)) || ((pixel_index2 >= 2332) && (pixel_index2 <= 2334)) || ((pixel_index2 >= 2341) && (pixel_index2 <= 2355)) || ((pixel_index2 >= 2374) && (pixel_index2 <= 2384)) || ((pixel_index2 >= 2392) && (pixel_index2 <= 2398)) || ((pixel_index2 >= 2428) && (pixel_index2 <= 2437)) || ((pixel_index2 >= 2443) && (pixel_index2 <= 2451)) || ((pixel_index2 >= 2470) && (pixel_index2 <= 2480)) || ((pixel_index2 >= 2487) && (pixel_index2 <= 2494)) || ((pixel_index2 >= 2526) && (pixel_index2 <= 2532)) || ((pixel_index2 >= 2540) && (pixel_index2 <= 2547)) || pixel_index2 == 2566 || ((pixel_index2 >= 2580) && (pixel_index2 <= 2588)) || ((pixel_index2 >= 2622) && (pixel_index2 <= 2626)) || pixel_index2 == 2636 || ((pixel_index2 >= 2639) && (pixel_index2 <= 2644)) || ((pixel_index2 >= 2647) && (pixel_index2 <= 2648)) || pixel_index2 == 2659 || ((pixel_index2 >= 2661) && (pixel_index2 <= 2662)) || ((pixel_index2 >= 2676) && (pixel_index2 <= 2684)) || ((pixel_index2 >= 2718) && (pixel_index2 <= 2721)) || pixel_index2 == 2732 || ((pixel_index2 >= 2735) && (pixel_index2 <= 2742)) || ((pixel_index2 >= 2756) && (pixel_index2 <= 2758)) || ((pixel_index2 >= 2772) && (pixel_index2 <= 2780)) || ((pixel_index2 >= 2814) && (pixel_index2 <= 2817)) || pixel_index2 == 2828 || ((pixel_index2 >= 2831) && (pixel_index2 <= 2838)) || ((pixel_index2 >= 2842) && (pixel_index2 <= 2848)) || ((pixel_index2 >= 2852) && (pixel_index2 <= 2859)) || ((pixel_index2 >= 2866) && (pixel_index2 <= 2876)) || ((pixel_index2 >= 2910) && (pixel_index2 <= 2913)) || pixel_index2 == 2924 || ((pixel_index2 >= 2927) && (pixel_index2 <= 2935)) || ((pixel_index2 >= 2938) && (pixel_index2 <= 2944)) || ((pixel_index2 >= 2947) && (pixel_index2 <= 2955)) || pixel_index2 == 2962 || ((pixel_index2 >= 2964) && (pixel_index2 <= 2972)) || ((pixel_index2 >= 3006) && (pixel_index2 <= 3013)) || ((pixel_index2 >= 3019) && (pixel_index2 <= 3021)) || ((pixel_index2 >= 3023) && (pixel_index2 <= 3032)) || ((pixel_index2 >= 3042) && (pixel_index2 <= 3051)) || ((pixel_index2 >= 3058) && (pixel_index2 <= 3060)) || pixel_index2 == 3063 || ((pixel_index2 >= 3065) && (pixel_index2 <= 3068)) || ((pixel_index2 >= 3102) && (pixel_index2 <= 3104)) || pixel_index2 == 3107 || ((pixel_index2 >= 3117) && (pixel_index2 <= 3123)) || ((pixel_index2 >= 3143) && (pixel_index2 <= 3147)) || ((pixel_index2 >= 3154) && (pixel_index2 <= 3155)) || pixel_index2 == 3159 || ((pixel_index2 >= 3161) && (pixel_index2 <= 3164)) || ((pixel_index2 >= 3198) && (pixel_index2 <= 3200)) || ((pixel_index2 >= 3202) && (pixel_index2 <= 3203)) || ((pixel_index2 >= 3213) && (pixel_index2 <= 3216)) || ((pixel_index2 >= 3218) && (pixel_index2 <= 3219)) || ((pixel_index2 >= 3239) && (pixel_index2 <= 3243)) || ((pixel_index2 >= 3250) && (pixel_index2 <= 3251)) || ((pixel_index2 >= 3255) && (pixel_index2 <= 3260)) || ((pixel_index2 >= 3292) && (pixel_index2 <= 3299)) || ((pixel_index2 >= 3309) && (pixel_index2 <= 3312)) || ((pixel_index2 >= 3314) && (pixel_index2 <= 3315)) || ((pixel_index2 >= 3335) && (pixel_index2 <= 3337)) || pixel_index2 == 3339 || ((pixel_index2 >= 3346) && (pixel_index2 <= 3347)) || ((pixel_index2 >= 3351) && (pixel_index2 <= 3352)) || ((pixel_index2 >= 3354) && (pixel_index2 <= 3358)) || ((pixel_index2 >= 3388) && (pixel_index2 <= 3393)) || pixel_index2 == 3395 || ((pixel_index2 >= 3405) && (pixel_index2 <= 3407)) || ((pixel_index2 >= 3409) && (pixel_index2 <= 3411)) || ((pixel_index2 >= 3431) && (pixel_index2 <= 3432)) || ((pixel_index2 >= 3434) && (pixel_index2 <= 3435)) || ((pixel_index2 >= 3438) && (pixel_index2 <= 3443)) || ((pixel_index2 >= 3447) && (pixel_index2 <= 3448)) || ((pixel_index2 >= 3450) && (pixel_index2 <= 3454)) || ((pixel_index2 >= 3484) && (pixel_index2 <= 3487)) || pixel_index2 == 3489 || pixel_index2 == 3491 || ((pixel_index2 >= 3501) && (pixel_index2 <= 3502)) || ((pixel_index2 >= 3505) && (pixel_index2 <= 3507)) || ((pixel_index2 >= 3527) && (pixel_index2 <= 3531)) || ((pixel_index2 >= 3538) && (pixel_index2 <= 3539)) || ((pixel_index2 >= 3543) && (pixel_index2 <= 3544)) || ((pixel_index2 >= 3546) && (pixel_index2 <= 3550)) || ((pixel_index2 >= 3580) && (pixel_index2 <= 3587)) || ((pixel_index2 >= 3597) && (pixel_index2 <= 3603)) || ((pixel_index2 >= 3623) && (pixel_index2 <= 3628)) || ((pixel_index2 >= 3633) && (pixel_index2 <= 3635)) || ((pixel_index2 >= 3639) && (pixel_index2 <= 3646)) || ((pixel_index2 >= 4620) && (pixel_index2 <= 4692)) || ((pixel_index2 >= 4707) && (pixel_index2 <= 4796)) || ((pixel_index2 >= 4803) && (pixel_index2 <= 4812)) || ((pixel_index2 >= 4814) && (pixel_index2 <= 4817)) || ((pixel_index2 >= 4819) && (pixel_index2 <= 4820)) || ((pixel_index2 >= 4827) && (pixel_index2 <= 4829)) || ((pixel_index2 >= 4834) && (pixel_index2 <= 4835)) || ((pixel_index2 >= 4838) && (pixel_index2 <= 4839)) || ((pixel_index2 >= 4841) && (pixel_index2 <= 4843)) || ((pixel_index2 >= 4845) && (pixel_index2 <= 4846)) || ((pixel_index2 >= 4851) && (pixel_index2 <= 4861)) || ((pixel_index2 >= 4863) && (pixel_index2 <= 4865)) || ((pixel_index2 >= 4868) && (pixel_index2 <= 4869)) || ((pixel_index2 >= 4871) && (pixel_index2 <= 4873)) || ((pixel_index2 >= 4880) && (pixel_index2 <= 4882)) || ((pixel_index2 >= 4887) && (pixel_index2 <= 4892)) || ((pixel_index2 >= 4899) && (pixel_index2 <= 4907)) || ((pixel_index2 >= 4910) && (pixel_index2 <= 4912)) || pixel_index2 == 4915 || pixel_index2 == 4924 || pixel_index2 == 4931 || pixel_index2 == 4935 || pixel_index2 == 4938 || pixel_index2 == 4941 || ((pixel_index2 >= 4948) && (pixel_index2 <= 4956)) || ((pixel_index2 >= 4959) && (pixel_index2 <= 4961)) || pixel_index2 == 4965 || pixel_index2 == 4968 || pixel_index2 == 4977 || ((pixel_index2 >= 4984) && (pixel_index2 <= 4988)) || ((pixel_index2 >= 4994) && (pixel_index2 <= 5003)) || ((pixel_index2 >= 5006) && (pixel_index2 <= 5008)) || pixel_index2 == 5011 || pixel_index2 == 5020 || pixel_index2 == 5027 || pixel_index2 == 5034 || pixel_index2 == 5037 || ((pixel_index2 >= 5044) && (pixel_index2 <= 5052)) || ((pixel_index2 >= 5055) && (pixel_index2 <= 5057)) || pixel_index2 == 5064 || pixel_index2 == 5073 || ((pixel_index2 >= 5080) && (pixel_index2 <= 5085)) || ((pixel_index2 >= 5090) && (pixel_index2 <= 5099)) || ((pixel_index2 >= 5102) && (pixel_index2 <= 5104)) || pixel_index2 == 5107 || ((pixel_index2 >= 5111) && (pixel_index2 <= 5112)) || ((pixel_index2 >= 5116) && (pixel_index2 <= 5119)) || ((pixel_index2 >= 5123) && (pixel_index2 <= 5124)) || pixel_index2 == 5130 || ((pixel_index2 >= 5133) && (pixel_index2 <= 5136)) || ((pixel_index2 >= 5140) && (pixel_index2 <= 5148)) || ((pixel_index2 >= 5151) && (pixel_index2 <= 5154)) || pixel_index2 == 5160 || ((pixel_index2 >= 5164) && (pixel_index2 <= 5165)) || pixel_index2 == 5169 || ((pixel_index2 >= 5173) && (pixel_index2 <= 5181)) || ((pixel_index2 >= 5186) && (pixel_index2 <= 5195)) || ((pixel_index2 >= 5198) && (pixel_index2 <= 5200)) || pixel_index2 == 5203 || ((pixel_index2 >= 5206) && (pixel_index2 <= 5209)) || ((pixel_index2 >= 5212) && (pixel_index2 <= 5216)) || ((pixel_index2 >= 5219) && (pixel_index2 <= 5220)) || pixel_index2 == 5226 || ((pixel_index2 >= 5229) && (pixel_index2 <= 5233)) || ((pixel_index2 >= 5236) && (pixel_index2 <= 5244)) || ((pixel_index2 >= 5247) && (pixel_index2 <= 5250)) || pixel_index2 == 5256 || ((pixel_index2 >= 5259) && (pixel_index2 <= 5262)) || pixel_index2 == 5265 || ((pixel_index2 >= 5271) && (pixel_index2 <= 5277)) || ((pixel_index2 >= 5282) && (pixel_index2 <= 5291)) || ((pixel_index2 >= 5294) && (pixel_index2 <= 5296)) || pixel_index2 == 5299 || ((pixel_index2 >= 5302) && (pixel_index2 <= 5305)) || ((pixel_index2 >= 5308) && (pixel_index2 <= 5312)) || pixel_index2 == 5315 || pixel_index2 == 5322 || ((pixel_index2 >= 5325) && (pixel_index2 <= 5329)) || ((pixel_index2 >= 5332) && (pixel_index2 <= 5340)) || ((pixel_index2 >= 5343) && (pixel_index2 <= 5345)) || pixel_index2 == 5352 || ((pixel_index2 >= 5355) && (pixel_index2 <= 5358)) || pixel_index2 == 5361 || ((pixel_index2 >= 5368) && (pixel_index2 <= 5373)) || ((pixel_index2 >= 5378) && (pixel_index2 <= 5387)) || ((pixel_index2 >= 5390) && (pixel_index2 <= 5392)) || pixel_index2 == 5395 || ((pixel_index2 >= 5398) && (pixel_index2 <= 5401)) || ((pixel_index2 >= 5404) && (pixel_index2 <= 5408)) || pixel_index2 == 5411 || pixel_index2 == 5415 || pixel_index2 == 5418 || ((pixel_index2 >= 5421) && (pixel_index2 <= 5425)) || ((pixel_index2 >= 5428) && (pixel_index2 <= 5436)) || ((pixel_index2 >= 5439) && (pixel_index2 <= 5441)) || pixel_index2 == 5445 || pixel_index2 == 5448 || ((pixel_index2 >= 5451) && (pixel_index2 <= 5454)) || ((pixel_index2 >= 5457) && (pixel_index2 <= 5458)) || ((pixel_index2 >= 5464) && (pixel_index2 <= 5469)) || ((pixel_index2 >= 5474) && (pixel_index2 <= 5483)) || ((pixel_index2 >= 5486) && (pixel_index2 <= 5488)) || pixel_index2 == 5491 || ((pixel_index2 >= 5494) && (pixel_index2 <= 5497)) || ((pixel_index2 >= 5500) && (pixel_index2 <= 5503)) || pixel_index2 == 5507 || ((pixel_index2 >= 5510) && (pixel_index2 <= 5511)) || pixel_index2 == 5514 || ((pixel_index2 >= 5517) && (pixel_index2 <= 5520)) || ((pixel_index2 >= 5524) && (pixel_index2 <= 5532)) || ((pixel_index2 >= 5535) && (pixel_index2 <= 5537)) || ((pixel_index2 >= 5540) && (pixel_index2 <= 5541)) || pixel_index2 == 5544 || ((pixel_index2 >= 5548) && (pixel_index2 <= 5549)) || ((pixel_index2 >= 5553) && (pixel_index2 <= 5556)) || ((pixel_index2 >= 5560) && (pixel_index2 <= 5565)) || ((pixel_index2 >= 5570) && (pixel_index2 <= 5575)) || pixel_index2 == 5584 || pixel_index2 == 5587 || ((pixel_index2 >= 5590) && (pixel_index2 <= 5593)) || pixel_index2 == 5596 || pixel_index2 == 5603 || pixel_index2 == 5610 || pixel_index2 == 5613 || ((pixel_index2 >= 5620) && (pixel_index2 <= 5624)) || pixel_index2 == 5633 || pixel_index2 == 5640 || pixel_index2 == 5649 || ((pixel_index2 >= 5656) && (pixel_index2 <= 5661)) || ((pixel_index2 >= 5667) && (pixel_index2 <= 5671)) || pixel_index2 == 5680 || pixel_index2 == 5683 || ((pixel_index2 >= 5686) && (pixel_index2 <= 5689)) || pixel_index2 == 5692 || pixel_index2 == 5699 || pixel_index2 == 5706 || pixel_index2 == 5709 || ((pixel_index2 >= 5716) && (pixel_index2 <= 5720)) || pixel_index2 == 5729 || pixel_index2 == 5736 || pixel_index2 == 5745 || ((pixel_index2 >= 5752) && (pixel_index2 <= 5756)) || ((pixel_index2 >= 5763) && (pixel_index2 <= 5768)) || ((pixel_index2 >= 5775) && (pixel_index2 <= 5776)) || ((pixel_index2 >= 5778) && (pixel_index2 <= 5780)) || ((pixel_index2 >= 5782) && (pixel_index2 <= 5785)) || ((pixel_index2 >= 5787) && (pixel_index2 <= 5789)) || ((pixel_index2 >= 5794) && (pixel_index2 <= 5796)) || ((pixel_index2 >= 5801) && (pixel_index2 <= 5802)) || ((pixel_index2 >= 5804) && (pixel_index2 <= 5806)) || ((pixel_index2 >= 5811) && (pixel_index2 <= 5817)) || ((pixel_index2 >= 5824) && (pixel_index2 <= 5826)) || ((pixel_index2 >= 5831) && (pixel_index2 <= 5833)) || ((pixel_index2 >= 5840) && (pixel_index2 <= 5842)) || ((pixel_index2 >= 5847) && (pixel_index2 <= 5852)) || (pixel_index2 >= 5868) && (pixel_index2 <= 5940)) oled_data2 = 16'b0000000000001010;
                    else if (((pixel_index2 >= 125) && (pixel_index2 <= 129)) || pixel_index2 == 221 || pixel_index2 == 225 || pixel_index2 == 317 || pixel_index2 == 321 || pixel_index2 == 413 || pixel_index2 == 417 || pixel_index2 == 509 || pixel_index2 == 513 || pixel_index2 == 605 || pixel_index2 == 609 || pixel_index2 == 701 || pixel_index2 == 705 || ((pixel_index2 >= 797) && (pixel_index2 <= 801)) || pixel_index2 == 1155 || ((pixel_index2 >= 1159) && (pixel_index2 <= 1161)) || pixel_index2 == 1163 || ((pixel_index2 >= 1165) && (pixel_index2 <= 1166)) || pixel_index2 == 1168 || ((pixel_index2 >= 1170) && (pixel_index2 <= 1171)) || pixel_index2 == 1173 || ((pixel_index2 >= 1175) && (pixel_index2 <= 1176)) || pixel_index2 == 1178 || pixel_index2 == 1254 || ((pixel_index2 >= 1256) && (pixel_index2 <= 1257)) || pixel_index2 == 1259 || ((pixel_index2 >= 1261) && (pixel_index2 <= 1262)) || ((pixel_index2 >= 1264) && (pixel_index2 <= 1267)) || ((pixel_index2 >= 1270) && (pixel_index2 <= 1272)) || pixel_index2 == 1350 || ((pixel_index2 >= 1352) && (pixel_index2 <= 1353)) || pixel_index2 == 1355 || ((pixel_index2 >= 1357) && (pixel_index2 <= 1358)) || pixel_index2 == 1360 || ((pixel_index2 >= 1362) && (pixel_index2 <= 1363)) || pixel_index2 == 1365 || ((pixel_index2 >= 1367) && (pixel_index2 <= 1368)) || ((pixel_index2 >= 1447) && (pixel_index2 <= 1449)) || ((pixel_index2 >= 1451) && (pixel_index2 <= 1454)) || ((pixel_index2 >= 1456) && (pixel_index2 <= 1459)) || ((pixel_index2 >= 1461) && (pixel_index2 <= 1464)) || pixel_index2 == 1466) oled_data2 = 16'b1010001010010100;
                    else if (((pixel_index2 >= 185) && (pixel_index2 <= 189)) || pixel_index2 == 281 || pixel_index2 == 285 || pixel_index2 == 377 || pixel_index2 == 381 || pixel_index2 == 473 || pixel_index2 == 477 || pixel_index2 == 569 || pixel_index2 == 573 || pixel_index2 == 665 || pixel_index2 == 669 || pixel_index2 == 761 || pixel_index2 == 765 || ((pixel_index2 >= 857) && (pixel_index2 <= 861)) || ((pixel_index2 >= 4008) && (pixel_index2 <= 4009)) || ((pixel_index2 >= 4012) && (pixel_index2 <= 4015)) || ((pixel_index2 >= 4017) && (pixel_index2 <= 4020)) || ((pixel_index2 >= 4022) && (pixel_index2 <= 4025)) || pixel_index2 == 4027 || ((pixel_index2 >= 4029) && (pixel_index2 <= 4030)) || ((pixel_index2 >= 4104) && (pixel_index2 <= 4105)) || ((pixel_index2 >= 4110) && (pixel_index2 <= 4111)) || ((pixel_index2 >= 4113) && (pixel_index2 <= 4114)) || ((pixel_index2 >= 4120) && (pixel_index2 <= 4121)) || ((pixel_index2 >= 4124) && (pixel_index2 <= 4126)) || ((pixel_index2 >= 4200) && (pixel_index2 <= 4201)) || ((pixel_index2 >= 4204) && (pixel_index2 <= 4205)) || pixel_index2 == 4207 || ((pixel_index2 >= 4210) && (pixel_index2 <= 4212)) || ((pixel_index2 >= 4214) && (pixel_index2 <= 4215)) || pixel_index2 == 4217 || pixel_index2 == 4219 || ((pixel_index2 >= 4221) && (pixel_index2 <= 4222)) || ((pixel_index2 >= 4295) && (pixel_index2 <= 4298)) || ((pixel_index2 >= 4300) && (pixel_index2 <= 4303)) || ((pixel_index2 >= 4305) && (pixel_index2 <= 4307)) || ((pixel_index2 >= 4310) && (pixel_index2 <= 4313)) || (pixel_index2 >= 4315) && (pixel_index2 <= 4318)) oled_data2 = 16'b0101011110010100;
                    else if (pixel_index2 == 319 || pixel_index2 == 323 || pixel_index2 == 327 || pixel_index2 == 347 || pixel_index2 == 351 || pixel_index2 == 355 || pixel_index2 == 415 || pixel_index2 == 419 || pixel_index2 == 423 || pixel_index2 == 443 || pixel_index2 == 447 || pixel_index2 == 451 || pixel_index2 == 3253 || pixel_index2 == 3349) oled_data2 = 16'b0000010100000000;
                    else if (pixel_index2 == 523 || pixel_index2 == 527 || pixel_index2 == 531 || pixel_index2 == 535 || pixel_index2 == 551 || pixel_index2 == 555 || pixel_index2 == 559 || pixel_index2 == 563 || pixel_index2 == 567 || pixel_index2 == 571 || pixel_index2 == 619 || pixel_index2 == 623 || pixel_index2 == 627 || pixel_index2 == 631 || pixel_index2 == 647 || pixel_index2 == 651 || pixel_index2 == 655 || pixel_index2 == 659 || pixel_index2 == 663 || pixel_index2 == 667 || pixel_index2 == 3488) oled_data2 = 16'b1010000000000000;
                    else if (pixel_index2 == 1086 || pixel_index2 == 1098 || pixel_index2 == 1102 || pixel_index2 == 1106 || pixel_index2 == 1110 || pixel_index2 == 1126 || pixel_index2 == 1130 || pixel_index2 == 1134 || pixel_index2 == 1138 || pixel_index2 == 1142 || pixel_index2 == 1146) oled_data2 = 16'b0000001010000000;
                    else if (pixel_index2 == 1090 || pixel_index2 == 1094 || pixel_index2 == 1114 || pixel_index2 == 1118 || pixel_index2 == 1122) oled_data2 = 16'b1111011110001010;
                    else if (((pixel_index2 >= 1281) && (pixel_index2 <= 1282)) || pixel_index2 == 1292 || pixel_index2 == 1295 || ((pixel_index2 >= 1297) && (pixel_index2 <= 1299)) || pixel_index2 == 1302 || ((pixel_index2 >= 1304) && (pixel_index2 <= 1305)) || pixel_index2 == 1307 || pixel_index2 == 1309 || pixel_index2 == 1311 || pixel_index2 == 1313 || pixel_index2 == 1377 || ((pixel_index2 >= 1392) && (pixel_index2 <= 1395)) || ((pixel_index2 >= 1397) && (pixel_index2 <= 1399)) || pixel_index2 == 1401 || ((pixel_index2 >= 1403) && (pixel_index2 <= 1404)) || pixel_index2 == 1406 || pixel_index2 == 1409 || ((pixel_index2 >= 1487) && (pixel_index2 <= 1488)) || pixel_index2 == 1490 || pixel_index2 == 1493 || pixel_index2 == 1495 || pixel_index2 == 1497 || ((pixel_index2 >= 1499) && (pixel_index2 <= 1500)) || ((pixel_index2 >= 1502) && (pixel_index2 <= 1503)) || pixel_index2 == 1505 || pixel_index2 == 1697 || pixel_index2 == 1776 || ((pixel_index2 >= 1790) && (pixel_index2 <= 1791)) || pixel_index2 == 1793 || pixel_index2 == 1817 || pixel_index2 == 1871 || pixel_index2 == 1914 || pixel_index2 == 1974 || ((pixel_index2 >= 1989) && (pixel_index2 <= 1990)) || pixel_index2 == 1992 || pixel_index2 == 1995 || ((pixel_index2 >= 1997) && (pixel_index2 <= 1999)) || ((pixel_index2 >= 2009) && (pixel_index2 <= 2010)) || pixel_index2 == 2047 || ((pixel_index2 >= 2070) && (pixel_index2 <= 2071)) || pixel_index2 == 2083 || ((pixel_index2 >= 2086) && (pixel_index2 <= 2088)) || pixel_index2 == 2090 || pixel_index2 == 2094 || pixel_index2 == 2106 || pixel_index2 == 2141 || pixel_index2 == 2143 || ((pixel_index2 >= 2155) && (pixel_index2 <= 2156)) || pixel_index2 == 2179 || ((pixel_index2 >= 2185) && (pixel_index2 <= 2187)) || pixel_index2 == 2189 || pixel_index2 == 2240 || pixel_index2 == 2243 || pixel_index2 == 2251 || pixel_index2 == 2336 || pixel_index2 == 2338 || pixel_index2 == 2340 || pixel_index2 == 2548 || ((pixel_index2 >= 2550) && (pixel_index2 <= 2551)) || ((pixel_index2 >= 2562) && (pixel_index2 <= 2563)) || ((pixel_index2 >= 2567) && (pixel_index2 <= 2579)) || ((pixel_index2 >= 2645) && (pixel_index2 <= 2646)) || pixel_index2 == 2658 || pixel_index2 == 2660 || ((pixel_index2 >= 2663) && (pixel_index2 <= 2675)) || ((pixel_index2 >= 2759) && (pixel_index2 <= 2771)) || ((pixel_index2 >= 2925) && (pixel_index2 <= 2926)) || pixel_index2 == 2937 || pixel_index2 == 2946 || pixel_index2 == 3022 || ((pixel_index2 >= 3105) && (pixel_index2 <= 3106)) || pixel_index2 == 3201 || pixel_index2 == 3217 || ((pixel_index2 >= 3230) && (pixel_index2 <= 3231)) || pixel_index2 == 3313 || pixel_index2 == 3324 || pixel_index2 == 3408 || ((pixel_index2 >= 3421) && (pixel_index2 <= 3422)) || ((pixel_index2 >= 3503) && (pixel_index2 <= 3504)) || ((pixel_index2 >= 3533) && (pixel_index2 <= 3536)) || pixel_index2 == 3629 || pixel_index2 == 3632) oled_data2 = 16'b1010010100010100;
                    else if (pixel_index2 == 1287 || pixel_index2 == 1289 || pixel_index2 == 1479 || pixel_index2 == 1481 || pixel_index2 == 1667 || pixel_index2 == 1669 || pixel_index2 == 1671 || pixel_index2 == 1673 || pixel_index2 == 1675 || pixel_index2 == 1677 || pixel_index2 == 1859 || pixel_index2 == 1861 || pixel_index2 == 1863 || pixel_index2 == 1865 || pixel_index2 == 1867 || pixel_index2 == 1869 || ((pixel_index2 >= 1879) && (pixel_index2 <= 1881)) || ((pixel_index2 >= 1889) && (pixel_index2 <= 1891)) || ((pixel_index2 >= 1975) && (pixel_index2 <= 1987)) || ((pixel_index2 >= 2002) && (pixel_index2 <= 2007)) || pixel_index2 == 2055 || pixel_index2 == 2057 || ((pixel_index2 >= 2072) && (pixel_index2 <= 2073)) || ((pixel_index2 >= 2081) && (pixel_index2 <= 2082)) || ((pixel_index2 >= 2097) && (pixel_index2 <= 2103)) || pixel_index2 == 2169 || pixel_index2 == 2177 || ((pixel_index2 >= 2193) && (pixel_index2 <= 2194)) || ((pixel_index2 >= 2198) && (pixel_index2 <= 2199)) || pixel_index2 == 2239 || ((pixel_index2 >= 2241) && (pixel_index2 <= 2242)) || pixel_index2 == 2244 || pixel_index2 == 2247 || pixel_index2 == 2249 || pixel_index2 == 2265 || pixel_index2 == 2273 || ((pixel_index2 >= 2289) && (pixel_index2 <= 2290)) || ((pixel_index2 >= 2294) && (pixel_index2 <= 2295)) || pixel_index2 == 2335 || pixel_index2 == 2337 || pixel_index2 == 2339 || ((pixel_index2 >= 2356) && (pixel_index2 <= 2361)) || ((pixel_index2 >= 2369) && (pixel_index2 <= 2373)) || ((pixel_index2 >= 2385) && (pixel_index2 <= 2391)) || ((pixel_index2 >= 2438) && (pixel_index2 <= 2442)) || ((pixel_index2 >= 2452) && (pixel_index2 <= 2457)) || ((pixel_index2 >= 2465) && (pixel_index2 <= 2469)) || ((pixel_index2 >= 2481) && (pixel_index2 <= 2486)) || pixel_index2 == 2533 || pixel_index2 == 2539 || pixel_index2 == 2549 || ((pixel_index2 >= 2552) && (pixel_index2 <= 2553)) || pixel_index2 == 2561 || ((pixel_index2 >= 2564) && (pixel_index2 <= 2565)) || ((pixel_index2 >= 2627) && (pixel_index2 <= 2629)) || pixel_index2 == 2635 || ((pixel_index2 >= 2637) && (pixel_index2 <= 2638)) || pixel_index2 == 2649 || pixel_index2 == 2657 || ((pixel_index2 >= 2722) && (pixel_index2 <= 2725)) || pixel_index2 == 2731 || ((pixel_index2 >= 2733) && (pixel_index2 <= 2734)) || ((pixel_index2 >= 2743) && (pixel_index2 <= 2755)) || ((pixel_index2 >= 2818) && (pixel_index2 <= 2821)) || pixel_index2 == 2827 || ((pixel_index2 >= 2829) && (pixel_index2 <= 2830)) || ((pixel_index2 >= 2839) && (pixel_index2 <= 2841)) || ((pixel_index2 >= 2849) && (pixel_index2 <= 2851)) || ((pixel_index2 >= 2914) && (pixel_index2 <= 2917)) || pixel_index2 == 2923 || pixel_index2 == 2936 || pixel_index2 == 2945 || pixel_index2 == 2963 || ((pixel_index2 >= 3014) && (pixel_index2 <= 3018)) || ((pixel_index2 >= 3061) && (pixel_index2 <= 3062)) || pixel_index2 == 3064 || ((pixel_index2 >= 3108) && (pixel_index2 <= 3116)) || pixel_index2 == 3160 || ((pixel_index2 >= 3204) && (pixel_index2 <= 3212)) || ((pixel_index2 >= 3300) && (pixel_index2 <= 3308)) || pixel_index2 == 3317 || ((pixel_index2 >= 3319) && (pixel_index2 <= 3320)) || ((pixel_index2 >= 3330) && (pixel_index2 <= 3331)) || pixel_index2 == 3333 || pixel_index2 == 3338 || ((pixel_index2 >= 3396) && (pixel_index2 <= 3404)) || pixel_index2 == 3433 || ((pixel_index2 >= 3436) && (pixel_index2 <= 3437)) || ((pixel_index2 >= 3492) && (pixel_index2 <= 3500)) || ((pixel_index2 >= 3588) && (pixel_index2 <= 3596)) || ((pixel_index2 >= 3684) && (pixel_index2 <= 3692)) || ((pixel_index2 >= 3724) && (pixel_index2 <= 3729)) || ((pixel_index2 >= 3820) && (pixel_index2 <= 3825)) || ((pixel_index2 >= 3893) && (pixel_index2 <= 3894)) || ((pixel_index2 >= 3897) && (pixel_index2 <= 3905)) || ((pixel_index2 >= 3908) && (pixel_index2 <= 3909)) || ((pixel_index2 >= 3989) && (pixel_index2 <= 3990)) || ((pixel_index2 >= 3994) && (pixel_index2 <= 4000)) || ((pixel_index2 >= 4004) && (pixel_index2 <= 4005)) || ((pixel_index2 >= 4085) && (pixel_index2 <= 4086)) || ((pixel_index2 >= 4090) && (pixel_index2 <= 4096)) || ((pixel_index2 >= 4100) && (pixel_index2 <= 4101)) || pixel_index2 == 4706 || pixel_index2 == 4797 || pixel_index2 == 5666 || pixel_index2 == 5757) oled_data2 = 16'b0101001010001010;
                    else if (pixel_index2 == 1296 || ((pixel_index2 >= 1300) && (pixel_index2 <= 1301)) || pixel_index2 == 1303 || pixel_index2 == 1306 || pixel_index2 == 1308 || pixel_index2 == 1310 || pixel_index2 == 1312 || pixel_index2 == 1391 || pixel_index2 == 1396 || pixel_index2 == 1400 || pixel_index2 == 1402 || pixel_index2 == 1405 || ((pixel_index2 >= 1407) && (pixel_index2 <= 1408)) || pixel_index2 == 1489 || ((pixel_index2 >= 1491) && (pixel_index2 <= 1492)) || pixel_index2 == 1494 || pixel_index2 == 1496 || pixel_index2 == 1498 || pixel_index2 == 1501 || pixel_index2 == 1504 || pixel_index2 == 3353 || pixel_index2 == 3449 || pixel_index2 == 3545) oled_data2 = 16'b0101001010010100;
                    else if (pixel_index2 == 1319 || ((pixel_index2 >= 1322) && (pixel_index2 <= 1324)) || pixel_index2 == 1327 || pixel_index2 == 1329 || pixel_index2 == 1332 || pixel_index2 == 1415 || pixel_index2 == 1418 || pixel_index2 == 1423 || pixel_index2 == 1425 || pixel_index2 == 1428 || ((pixel_index2 >= 1509) && (pixel_index2 <= 1511)) || ((pixel_index2 >= 1514) && (pixel_index2 <= 1516)) || ((pixel_index2 >= 1519) && (pixel_index2 <= 1521)) || pixel_index2 == 1524 || pixel_index2 == 1612 || pixel_index2 == 1620 || ((pixel_index2 >= 1706) && (pixel_index2 <= 1708)) || pixel_index2 == 1716) oled_data2 = 16'b1010000000001010;
                    else if (((pixel_index2 >= 1570) && (pixel_index2 <= 1574)) || pixel_index2 == 1666 || pixel_index2 == 1670 || pixel_index2 == 1762 || pixel_index2 == 1766 || pixel_index2 == 1858 || pixel_index2 == 1862 || ((pixel_index2 >= 1954) && (pixel_index2 <= 1958)) || pixel_index2 == 2213 || pixel_index2 == 2216 || ((pixel_index2 >= 2219) && (pixel_index2 <= 2221)) || pixel_index2 == 2223 || pixel_index2 == 2226 || ((pixel_index2 >= 2228) && (pixel_index2 <= 2230)) || pixel_index2 == 2310 || pixel_index2 == 2312 || pixel_index2 == 2314 || pixel_index2 == 2319 || pixel_index2 == 2322 || pixel_index2 == 2325 || pixel_index2 == 2329 || ((pixel_index2 >= 2406) && (pixel_index2 <= 2408)) || ((pixel_index2 >= 2411) && (pixel_index2 <= 2412)) || ((pixel_index2 >= 2415) && (pixel_index2 <= 2416)) || pixel_index2 == 2418 || pixel_index2 == 2421 || pixel_index2 == 2424 || pixel_index2 == 2501 || pixel_index2 == 2504 || pixel_index2 == 2509 || pixel_index2 == 2511 || ((pixel_index2 >= 2513) && (pixel_index2 <= 2514)) || pixel_index2 == 2517 || pixel_index2 == 2521 || ((pixel_index2 >= 2598) && (pixel_index2 <= 2600)) || ((pixel_index2 >= 2602) && (pixel_index2 <= 2604)) || pixel_index2 == 2607 || pixel_index2 == 2610 || (pixel_index2 >= 2612) && (pixel_index2 <= 2614)) oled_data2 = 16'b1010011110001010;
                    else if (pixel_index2 == 3229 || (pixel_index2 >= 3325) && (pixel_index2 <= 3326)) oled_data2 = 16'b0101010100001010;
                    else if (pixel_index2 == 3394 || pixel_index2 == 3490) oled_data2 = 16'b0000000000010100;
                    else if (pixel_index2 == 3532 || pixel_index2 == 3537) oled_data2 = 16'b0101000000000000;
                    else if (((pixel_index2 >= 4423) && (pixel_index2 <= 4505)) || ((pixel_index2 >= 4513) && (pixel_index2 <= 4518)) || (pixel_index2 >= 4602) && (pixel_index2 <= 4606)) oled_data2 = 16'b0000001010011110;
                    else if (((pixel_index2 >= 4519) && (pixel_index2 <= 4601)) || ((pixel_index2 >= 4609) && (pixel_index2 <= 4619)) || ((pixel_index2 >= 4693) && (pixel_index2 <= 4702)) || pixel_index2 == 4705 || pixel_index2 == 4798 || pixel_index2 == 4801 || pixel_index2 == 4894 || ((pixel_index2 >= 4897) && (pixel_index2 <= 4898)) || ((pixel_index2 >= 4989) && (pixel_index2 <= 4990)) || pixel_index2 == 4993 || pixel_index2 == 5086 || pixel_index2 == 5089 || pixel_index2 == 5182 || pixel_index2 == 5185 || pixel_index2 == 5278 || pixel_index2 == 5281 || pixel_index2 == 5374 || pixel_index2 == 5377 || pixel_index2 == 5470 || pixel_index2 == 5473 || pixel_index2 == 5566 || pixel_index2 == 5569 || pixel_index2 == 5662 || pixel_index2 == 5665 || pixel_index2 == 5758 || pixel_index2 == 5761 || pixel_index2 == 5854 || ((pixel_index2 >= 5857) && (pixel_index2 <= 5867)) || ((pixel_index2 >= 5941) && (pixel_index2 <= 5950)) || (pixel_index2 >= 5959) && (pixel_index2 <= 6041)) oled_data2 = 16'b0000001010010100;
                    else if (pixel_index2 == 4813 || pixel_index2 == 4818 || ((pixel_index2 >= 4821) && (pixel_index2 <= 4826)) || ((pixel_index2 >= 4830) && (pixel_index2 <= 4833)) || ((pixel_index2 >= 4836) && (pixel_index2 <= 4837)) || pixel_index2 == 4840 || pixel_index2 == 4844 || ((pixel_index2 >= 4847) && (pixel_index2 <= 4850)) || pixel_index2 == 4862 || ((pixel_index2 >= 4866) && (pixel_index2 <= 4867)) || pixel_index2 == 4870 || ((pixel_index2 >= 4874) && (pixel_index2 <= 4879)) || ((pixel_index2 >= 4883) && (pixel_index2 <= 4886)) || pixel_index2 == 4908 || pixel_index2 == 4913 || pixel_index2 == 4916 || pixel_index2 == 4923 || pixel_index2 == 4925 || pixel_index2 == 4930 || pixel_index2 == 4934 || pixel_index2 == 4937 || pixel_index2 == 4939 || pixel_index2 == 4942 || pixel_index2 == 4947 || pixel_index2 == 4957 || pixel_index2 == 4964 || pixel_index2 == 4967 || pixel_index2 == 4969 || pixel_index2 == 4976 || pixel_index2 == 4978 || pixel_index2 == 4983 || pixel_index2 == 5031 || pixel_index2 == 5061 || pixel_index2 == 5221 || pixel_index2 == 5251 || ((pixel_index2 >= 5268) && (pixel_index2 <= 5270)) || pixel_index2 == 5316 || pixel_index2 == 5346 || pixel_index2 == 5367 || pixel_index2 == 5504 || pixel_index2 == 5521 || pixel_index2 == 5547 || pixel_index2 == 5550 || pixel_index2 == 5557 || ((pixel_index2 >= 5576) && (pixel_index2 <= 5579)) || ((pixel_index2 >= 5582) && (pixel_index2 <= 5583)) || ((pixel_index2 >= 5597) && (pixel_index2 <= 5599)) || ((pixel_index2 >= 5606) && (pixel_index2 <= 5607)) || ((pixel_index2 >= 5614) && (pixel_index2 <= 5616)) || ((pixel_index2 >= 5625) && (pixel_index2 <= 5628)) || ((pixel_index2 >= 5631) && (pixel_index2 <= 5632)) || ((pixel_index2 >= 5636) && (pixel_index2 <= 5637)) || ((pixel_index2 >= 5644) && (pixel_index2 <= 5645)) || (pixel_index2 >= 5650) && (pixel_index2 <= 5652)) oled_data2 = 16'b0101001010000000;
                    else if (pixel_index2 == 4909 || pixel_index2 == 4914 || ((pixel_index2 >= 4917) && (pixel_index2 <= 4922)) || ((pixel_index2 >= 4926) && (pixel_index2 <= 4929)) || ((pixel_index2 >= 4932) && (pixel_index2 <= 4933)) || pixel_index2 == 4936 || pixel_index2 == 4940 || ((pixel_index2 >= 4943) && (pixel_index2 <= 4946)) || pixel_index2 == 4958 || ((pixel_index2 >= 4962) && (pixel_index2 <= 4963)) || pixel_index2 == 4966 || ((pixel_index2 >= 4970) && (pixel_index2 <= 4975)) || ((pixel_index2 >= 4979) && (pixel_index2 <= 4982)) || ((pixel_index2 >= 5004) && (pixel_index2 <= 5005)) || ((pixel_index2 >= 5009) && (pixel_index2 <= 5010)) || ((pixel_index2 >= 5012) && (pixel_index2 <= 5019)) || ((pixel_index2 >= 5021) && (pixel_index2 <= 5026)) || ((pixel_index2 >= 5028) && (pixel_index2 <= 5030)) || ((pixel_index2 >= 5032) && (pixel_index2 <= 5033)) || ((pixel_index2 >= 5035) && (pixel_index2 <= 5036)) || ((pixel_index2 >= 5038) && (pixel_index2 <= 5043)) || ((pixel_index2 >= 5053) && (pixel_index2 <= 5054)) || ((pixel_index2 >= 5058) && (pixel_index2 <= 5060)) || ((pixel_index2 >= 5062) && (pixel_index2 <= 5063)) || ((pixel_index2 >= 5065) && (pixel_index2 <= 5072)) || ((pixel_index2 >= 5074) && (pixel_index2 <= 5079)) || ((pixel_index2 >= 5100) && (pixel_index2 <= 5101)) || ((pixel_index2 >= 5105) && (pixel_index2 <= 5106)) || ((pixel_index2 >= 5108) && (pixel_index2 <= 5110)) || ((pixel_index2 >= 5113) && (pixel_index2 <= 5115)) || ((pixel_index2 >= 5120) && (pixel_index2 <= 5122)) || ((pixel_index2 >= 5125) && (pixel_index2 <= 5129)) || ((pixel_index2 >= 5131) && (pixel_index2 <= 5132)) || ((pixel_index2 >= 5137) && (pixel_index2 <= 5139)) || ((pixel_index2 >= 5149) && (pixel_index2 <= 5150)) || ((pixel_index2 >= 5155) && (pixel_index2 <= 5159)) || ((pixel_index2 >= 5161) && (pixel_index2 <= 5163)) || ((pixel_index2 >= 5166) && (pixel_index2 <= 5168)) || ((pixel_index2 >= 5170) && (pixel_index2 <= 5172)) || ((pixel_index2 >= 5196) && (pixel_index2 <= 5197)) || ((pixel_index2 >= 5201) && (pixel_index2 <= 5202)) || ((pixel_index2 >= 5204) && (pixel_index2 <= 5205)) || ((pixel_index2 >= 5210) && (pixel_index2 <= 5211)) || ((pixel_index2 >= 5217) && (pixel_index2 <= 5218)) || ((pixel_index2 >= 5222) && (pixel_index2 <= 5225)) || ((pixel_index2 >= 5227) && (pixel_index2 <= 5228)) || ((pixel_index2 >= 5234) && (pixel_index2 <= 5235)) || ((pixel_index2 >= 5245) && (pixel_index2 <= 5246)) || ((pixel_index2 >= 5252) && (pixel_index2 <= 5255)) || ((pixel_index2 >= 5257) && (pixel_index2 <= 5258)) || ((pixel_index2 >= 5263) && (pixel_index2 <= 5264)) || ((pixel_index2 >= 5266) && (pixel_index2 <= 5267)) || ((pixel_index2 >= 5292) && (pixel_index2 <= 5293)) || ((pixel_index2 >= 5297) && (pixel_index2 <= 5298)) || ((pixel_index2 >= 5300) && (pixel_index2 <= 5301)) || ((pixel_index2 >= 5306) && (pixel_index2 <= 5307)) || ((pixel_index2 >= 5313) && (pixel_index2 <= 5314)) || ((pixel_index2 >= 5317) && (pixel_index2 <= 5321)) || ((pixel_index2 >= 5323) && (pixel_index2 <= 5324)) || ((pixel_index2 >= 5330) && (pixel_index2 <= 5331)) || ((pixel_index2 >= 5341) && (pixel_index2 <= 5342)) || ((pixel_index2 >= 5347) && (pixel_index2 <= 5351)) || ((pixel_index2 >= 5353) && (pixel_index2 <= 5354)) || ((pixel_index2 >= 5359) && (pixel_index2 <= 5360)) || ((pixel_index2 >= 5362) && (pixel_index2 <= 5366)) || ((pixel_index2 >= 5388) && (pixel_index2 <= 5389)) || ((pixel_index2 >= 5393) && (pixel_index2 <= 5394)) || ((pixel_index2 >= 5396) && (pixel_index2 <= 5397)) || ((pixel_index2 >= 5402) && (pixel_index2 <= 5403)) || ((pixel_index2 >= 5409) && (pixel_index2 <= 5410)) || ((pixel_index2 >= 5412) && (pixel_index2 <= 5414)) || ((pixel_index2 >= 5416) && (pixel_index2 <= 5417)) || ((pixel_index2 >= 5419) && (pixel_index2 <= 5420)) || ((pixel_index2 >= 5426) && (pixel_index2 <= 5427)) || ((pixel_index2 >= 5437) && (pixel_index2 <= 5438)) || ((pixel_index2 >= 5442) && (pixel_index2 <= 5444)) || ((pixel_index2 >= 5446) && (pixel_index2 <= 5447)) || ((pixel_index2 >= 5449) && (pixel_index2 <= 5450)) || ((pixel_index2 >= 5455) && (pixel_index2 <= 5456)) || ((pixel_index2 >= 5459) && (pixel_index2 <= 5463)) || ((pixel_index2 >= 5484) && (pixel_index2 <= 5485)) || ((pixel_index2 >= 5489) && (pixel_index2 <= 5490)) || ((pixel_index2 >= 5492) && (pixel_index2 <= 5493)) || ((pixel_index2 >= 5498) && (pixel_index2 <= 5499)) || ((pixel_index2 >= 5505) && (pixel_index2 <= 5506)) || ((pixel_index2 >= 5508) && (pixel_index2 <= 5509)) || ((pixel_index2 >= 5512) && (pixel_index2 <= 5513)) || ((pixel_index2 >= 5515) && (pixel_index2 <= 5516)) || ((pixel_index2 >= 5522) && (pixel_index2 <= 5523)) || ((pixel_index2 >= 5533) && (pixel_index2 <= 5534)) || ((pixel_index2 >= 5538) && (pixel_index2 <= 5539)) || ((pixel_index2 >= 5542) && (pixel_index2 <= 5543)) || ((pixel_index2 >= 5545) && (pixel_index2 <= 5546)) || ((pixel_index2 >= 5551) && (pixel_index2 <= 5552)) || ((pixel_index2 >= 5558) && (pixel_index2 <= 5559)) || ((pixel_index2 >= 5580) && (pixel_index2 <= 5581)) || ((pixel_index2 >= 5585) && (pixel_index2 <= 5586)) || ((pixel_index2 >= 5588) && (pixel_index2 <= 5589)) || ((pixel_index2 >= 5594) && (pixel_index2 <= 5595)) || ((pixel_index2 >= 5600) && (pixel_index2 <= 5602)) || ((pixel_index2 >= 5604) && (pixel_index2 <= 5605)) || ((pixel_index2 >= 5608) && (pixel_index2 <= 5609)) || ((pixel_index2 >= 5611) && (pixel_index2 <= 5612)) || ((pixel_index2 >= 5617) && (pixel_index2 <= 5619)) || ((pixel_index2 >= 5629) && (pixel_index2 <= 5630)) || ((pixel_index2 >= 5634) && (pixel_index2 <= 5635)) || ((pixel_index2 >= 5638) && (pixel_index2 <= 5639)) || ((pixel_index2 >= 5641) && (pixel_index2 <= 5643)) || ((pixel_index2 >= 5646) && (pixel_index2 <= 5648)) || ((pixel_index2 >= 5653) && (pixel_index2 <= 5655)) || ((pixel_index2 >= 5672) && (pixel_index2 <= 5679)) || ((pixel_index2 >= 5681) && (pixel_index2 <= 5682)) || ((pixel_index2 >= 5684) && (pixel_index2 <= 5685)) || ((pixel_index2 >= 5690) && (pixel_index2 <= 5691)) || ((pixel_index2 >= 5693) && (pixel_index2 <= 5698)) || ((pixel_index2 >= 5700) && (pixel_index2 <= 5705)) || ((pixel_index2 >= 5707) && (pixel_index2 <= 5708)) || ((pixel_index2 >= 5710) && (pixel_index2 <= 5715)) || ((pixel_index2 >= 5721) && (pixel_index2 <= 5728)) || ((pixel_index2 >= 5730) && (pixel_index2 <= 5735)) || ((pixel_index2 >= 5737) && (pixel_index2 <= 5744)) || ((pixel_index2 >= 5746) && (pixel_index2 <= 5751)) || ((pixel_index2 >= 5769) && (pixel_index2 <= 5774)) || pixel_index2 == 5777 || pixel_index2 == 5781 || pixel_index2 == 5786 || ((pixel_index2 >= 5790) && (pixel_index2 <= 5793)) || ((pixel_index2 >= 5797) && (pixel_index2 <= 5800)) || pixel_index2 == 5803 || ((pixel_index2 >= 5807) && (pixel_index2 <= 5810)) || ((pixel_index2 >= 5818) && (pixel_index2 <= 5823)) || ((pixel_index2 >= 5827) && (pixel_index2 <= 5830)) || ((pixel_index2 >= 5834) && (pixel_index2 <= 5839)) || (pixel_index2 >= 5843) && (pixel_index2 <= 5846)) oled_data2 = 16'b1111010100010100;
                    else oled_data2 = 0;
                end
                6: begin
                    if (pixel_index2 == 97 || pixel_index2 == 99 || pixel_index2 == 101 || ((pixel_index2 >= 103) && (pixel_index2 <= 104)) || ((pixel_index2 >= 106) && (pixel_index2 <= 109)) || pixel_index2 == 111 || ((pixel_index2 >= 113) && (pixel_index2 <= 114)) || ((pixel_index2 >= 118) && (pixel_index2 <= 120)) || ((pixel_index2 >= 129) && (pixel_index2 <= 165)) || pixel_index2 == 195 || pixel_index2 == 197 || ((pixel_index2 >= 199) && (pixel_index2 <= 200)) || pixel_index2 == 202 || ((pixel_index2 >= 204) && (pixel_index2 <= 205)) || pixel_index2 == 207 || ((pixel_index2 >= 209) && (pixel_index2 <= 210)) || pixel_index2 == 213 || pixel_index2 == 225 || pixel_index2 == 261 || pixel_index2 == 289 || ((pixel_index2 >= 291) && (pixel_index2 <= 296)) || pixel_index2 == 298 || ((pixel_index2 >= 300) && (pixel_index2 <= 301)) || pixel_index2 == 303 || ((pixel_index2 >= 305) && (pixel_index2 <= 306)) || ((pixel_index2 >= 310) && (pixel_index2 <= 312)) || pixel_index2 == 321 || pixel_index2 == 357 || pixel_index2 == 385 || ((pixel_index2 >= 387) && (pixel_index2 <= 392)) || pixel_index2 == 394 || ((pixel_index2 >= 396) && (pixel_index2 <= 397)) || ((pixel_index2 >= 399) && (pixel_index2 <= 402)) || pixel_index2 == 408 || pixel_index2 == 417 || pixel_index2 == 453 || ((pixel_index2 >= 501) && (pixel_index2 <= 504)) || pixel_index2 == 513 || pixel_index2 == 549 || pixel_index2 == 609 || pixel_index2 == 645 || ((pixel_index2 >= 674) && (pixel_index2 <= 675)) || ((pixel_index2 >= 678) && (pixel_index2 <= 681)) || ((pixel_index2 >= 685) && (pixel_index2 <= 686)) || pixel_index2 == 688 || ((pixel_index2 >= 690) && (pixel_index2 <= 691)) || ((pixel_index2 >= 693) && (pixel_index2 <= 696)) || pixel_index2 == 698 || pixel_index2 == 705 || pixel_index2 == 741 || ((pixel_index2 >= 770) && (pixel_index2 <= 771)) || pixel_index2 == 774 || ((pixel_index2 >= 776) && (pixel_index2 <= 777)) || ((pixel_index2 >= 779) && (pixel_index2 <= 782)) || pixel_index2 == 784 || ((pixel_index2 >= 786) && (pixel_index2 <= 787)) || ((pixel_index2 >= 790) && (pixel_index2 <= 791)) || ((pixel_index2 >= 801) && (pixel_index2 <= 837)) || ((pixel_index2 >= 866) && (pixel_index2 <= 867)) || pixel_index2 == 870 || ((pixel_index2 >= 872) && (pixel_index2 <= 873)) || pixel_index2 == 875 || ((pixel_index2 >= 877) && (pixel_index2 <= 878)) || pixel_index2 == 880 || ((pixel_index2 >= 882) && (pixel_index2 <= 883)) || ((pixel_index2 >= 886) && (pixel_index2 <= 887)) || ((pixel_index2 >= 961) && (pixel_index2 <= 964)) || pixel_index2 == 966 || ((pixel_index2 >= 968) && (pixel_index2 <= 969)) || ((pixel_index2 >= 971) && (pixel_index2 <= 974)) || ((pixel_index2 >= 976) && (pixel_index2 <= 979)) || ((pixel_index2 >= 981) && (pixel_index2 <= 984)) || pixel_index2 == 986) oled_data2 = 16'b1111001010010100;
                    else if (((pixel_index2 >= 124) && (pixel_index2 <= 128)) || ((pixel_index2 >= 166) && (pixel_index2 <= 190)) || ((pixel_index2 >= 220) && (pixel_index2 <= 221)) || pixel_index2 == 229 || pixel_index2 == 233 || pixel_index2 == 237 || pixel_index2 == 241 || pixel_index2 == 245 || pixel_index2 == 249 || pixel_index2 == 253 || pixel_index2 == 257 || pixel_index2 == 265 || pixel_index2 == 269 || pixel_index2 == 273 || pixel_index2 == 277 || pixel_index2 == 281 || ((pixel_index2 >= 285) && (pixel_index2 <= 286)) || ((pixel_index2 >= 316) && (pixel_index2 <= 317)) || pixel_index2 == 325 || pixel_index2 == 329 || pixel_index2 == 333 || pixel_index2 == 337 || pixel_index2 == 341 || pixel_index2 == 345 || pixel_index2 == 349 || pixel_index2 == 353 || pixel_index2 == 361 || pixel_index2 == 365 || pixel_index2 == 369 || pixel_index2 == 373 || pixel_index2 == 377 || ((pixel_index2 >= 381) && (pixel_index2 <= 382)) || ((pixel_index2 >= 412) && (pixel_index2 <= 413)) || pixel_index2 == 421 || pixel_index2 == 425 || pixel_index2 == 429 || pixel_index2 == 433 || pixel_index2 == 437 || pixel_index2 == 441 || pixel_index2 == 445 || pixel_index2 == 449 || pixel_index2 == 457 || pixel_index2 == 461 || pixel_index2 == 465 || pixel_index2 == 469 || pixel_index2 == 473 || ((pixel_index2 >= 477) && (pixel_index2 <= 478)) || ((pixel_index2 >= 508) && (pixel_index2 <= 509)) || pixel_index2 == 517 || pixel_index2 == 521 || pixel_index2 == 525 || pixel_index2 == 529 || pixel_index2 == 533 || pixel_index2 == 537 || pixel_index2 == 541 || pixel_index2 == 545 || pixel_index2 == 553 || pixel_index2 == 557 || pixel_index2 == 561 || pixel_index2 == 565 || pixel_index2 == 569 || ((pixel_index2 >= 573) && (pixel_index2 <= 574)) || ((pixel_index2 >= 604) && (pixel_index2 <= 605)) || pixel_index2 == 613 || pixel_index2 == 617 || pixel_index2 == 621 || pixel_index2 == 625 || pixel_index2 == 629 || pixel_index2 == 633 || pixel_index2 == 637 || pixel_index2 == 641 || pixel_index2 == 649 || pixel_index2 == 653 || pixel_index2 == 657 || pixel_index2 == 661 || pixel_index2 == 665 || ((pixel_index2 >= 669) && (pixel_index2 <= 670)) || ((pixel_index2 >= 700) && (pixel_index2 <= 701)) || pixel_index2 == 709 || pixel_index2 == 713 || pixel_index2 == 717 || pixel_index2 == 721 || pixel_index2 == 725 || pixel_index2 == 729 || pixel_index2 == 733 || pixel_index2 == 737 || pixel_index2 == 745 || pixel_index2 == 749 || pixel_index2 == 753 || pixel_index2 == 757 || pixel_index2 == 761 || ((pixel_index2 >= 765) && (pixel_index2 <= 766)) || ((pixel_index2 >= 796) && (pixel_index2 <= 800)) || ((pixel_index2 >= 838) && (pixel_index2 <= 862)) || ((pixel_index2 >= 892) && (pixel_index2 <= 894)) || ((pixel_index2 >= 897) && (pixel_index2 <= 898)) || ((pixel_index2 >= 901) && (pixel_index2 <= 902)) || ((pixel_index2 >= 905) && (pixel_index2 <= 906)) || ((pixel_index2 >= 909) && (pixel_index2 <= 910)) || ((pixel_index2 >= 913) && (pixel_index2 <= 914)) || ((pixel_index2 >= 917) && (pixel_index2 <= 918)) || ((pixel_index2 >= 921) && (pixel_index2 <= 922)) || ((pixel_index2 >= 925) && (pixel_index2 <= 926)) || ((pixel_index2 >= 929) && (pixel_index2 <= 930)) || ((pixel_index2 >= 933) && (pixel_index2 <= 934)) || ((pixel_index2 >= 937) && (pixel_index2 <= 938)) || ((pixel_index2 >= 941) && (pixel_index2 <= 942)) || ((pixel_index2 >= 945) && (pixel_index2 <= 946)) || ((pixel_index2 >= 949) && (pixel_index2 <= 950)) || ((pixel_index2 >= 953) && (pixel_index2 <= 954)) || ((pixel_index2 >= 957) && (pixel_index2 <= 958)) || ((pixel_index2 >= 988) && (pixel_index2 <= 1054)) || ((pixel_index2 >= 1084) && (pixel_index2 <= 1085)) || ((pixel_index2 >= 1087) && (pixel_index2 <= 1089)) || ((pixel_index2 >= 1091) && (pixel_index2 <= 1093)) || ((pixel_index2 >= 1095) && (pixel_index2 <= 1097)) || ((pixel_index2 >= 1099) && (pixel_index2 <= 1101)) || ((pixel_index2 >= 1103) && (pixel_index2 <= 1105)) || ((pixel_index2 >= 1107) && (pixel_index2 <= 1109)) || ((pixel_index2 >= 1111) && (pixel_index2 <= 1113)) || ((pixel_index2 >= 1115) && (pixel_index2 <= 1117)) || ((pixel_index2 >= 1119) && (pixel_index2 <= 1121)) || ((pixel_index2 >= 1123) && (pixel_index2 <= 1125)) || ((pixel_index2 >= 1127) && (pixel_index2 <= 1129)) || ((pixel_index2 >= 1131) && (pixel_index2 <= 1133)) || ((pixel_index2 >= 1135) && (pixel_index2 <= 1137)) || ((pixel_index2 >= 1139) && (pixel_index2 <= 1141)) || ((pixel_index2 >= 1143) && (pixel_index2 <= 1145)) || ((pixel_index2 >= 1147) && (pixel_index2 <= 1150)) || ((pixel_index2 >= 1182) && (pixel_index2 <= 1189)) || ((pixel_index2 >= 1195) && (pixel_index2 <= 1219)) || ((pixel_index2 >= 1240) && (pixel_index2 <= 1244)) || ((pixel_index2 >= 1278) && (pixel_index2 <= 1280)) || ((pixel_index2 >= 1283) && (pixel_index2 <= 1285)) || pixel_index2 == 1291 || ((pixel_index2 >= 1293) && (pixel_index2 <= 1294)) || ((pixel_index2 >= 1314) && (pixel_index2 <= 1315)) || ((pixel_index2 >= 1336) && (pixel_index2 <= 1340)) || ((pixel_index2 >= 1374) && (pixel_index2 <= 1376)) || ((pixel_index2 >= 1378) && (pixel_index2 <= 1381)) || ((pixel_index2 >= 1387) && (pixel_index2 <= 1390)) || ((pixel_index2 >= 1410) && (pixel_index2 <= 1411)) || ((pixel_index2 >= 1432) && (pixel_index2 <= 1436)) || ((pixel_index2 >= 1470) && (pixel_index2 <= 1477)) || ((pixel_index2 >= 1483) && (pixel_index2 <= 1486)) || ((pixel_index2 >= 1506) && (pixel_index2 <= 1507)) || ((pixel_index2 >= 1528) && (pixel_index2 <= 1532)) || ((pixel_index2 >= 1566) && (pixel_index2 <= 1573)) || ((pixel_index2 >= 1579) && (pixel_index2 <= 1603)) || ((pixel_index2 >= 1624) && (pixel_index2 <= 1628)) || ((pixel_index2 >= 1662) && (pixel_index2 <= 1666)) || pixel_index2 == 1670 || pixel_index2 == 1674 || ((pixel_index2 >= 1678) && (pixel_index2 <= 1696)) || ((pixel_index2 >= 1698) && (pixel_index2 <= 1699)) || ((pixel_index2 >= 1720) && (pixel_index2 <= 1724)) || ((pixel_index2 >= 1758) && (pixel_index2 <= 1762)) || pixel_index2 == 1766 || pixel_index2 == 1770 || ((pixel_index2 >= 1774) && (pixel_index2 <= 1775)) || ((pixel_index2 >= 1777) && (pixel_index2 <= 1789)) || pixel_index2 == 1792 || ((pixel_index2 >= 1794) && (pixel_index2 <= 1795)) || pixel_index2 == 1816 || ((pixel_index2 >= 1818) && (pixel_index2 <= 1820)) || ((pixel_index2 >= 1854) && (pixel_index2 <= 1858)) || pixel_index2 == 1862 || pixel_index2 == 1866 || pixel_index2 == 1870 || ((pixel_index2 >= 1872) && (pixel_index2 <= 1878)) || ((pixel_index2 >= 1882) && (pixel_index2 <= 1888)) || ((pixel_index2 >= 1892) && (pixel_index2 <= 1913)) || ((pixel_index2 >= 1915) && (pixel_index2 <= 1916)) || ((pixel_index2 >= 1948) && (pixel_index2 <= 1973)) || pixel_index2 == 1988 || pixel_index2 == 1991 || ((pixel_index2 >= 1993) && (pixel_index2 <= 1994)) || pixel_index2 == 1996 || ((pixel_index2 >= 2000) && (pixel_index2 <= 2001)) || pixel_index2 == 2008 || ((pixel_index2 >= 2011) && (pixel_index2 <= 2014)) || ((pixel_index2 >= 2044) && (pixel_index2 <= 2046)) || ((pixel_index2 >= 2048) && (pixel_index2 <= 2054)) || ((pixel_index2 >= 2058) && (pixel_index2 <= 2069)) || ((pixel_index2 >= 2084) && (pixel_index2 <= 2085)) || pixel_index2 == 2089 || ((pixel_index2 >= 2091) && (pixel_index2 <= 2093)) || ((pixel_index2 >= 2095) && (pixel_index2 <= 2096)) || ((pixel_index2 >= 2104) && (pixel_index2 <= 2105)) || ((pixel_index2 >= 2107) && (pixel_index2 <= 2110)) || pixel_index2 == 2140 || pixel_index2 == 2142 || ((pixel_index2 >= 2144) && (pixel_index2 <= 2150)) || pixel_index2 == 2154 || ((pixel_index2 >= 2157) && (pixel_index2 <= 2168)) || pixel_index2 == 2178 || ((pixel_index2 >= 2180) && (pixel_index2 <= 2184)) || pixel_index2 == 2188 || ((pixel_index2 >= 2190) && (pixel_index2 <= 2192)) || ((pixel_index2 >= 2195) && (pixel_index2 <= 2197)) || ((pixel_index2 >= 2200) && (pixel_index2 <= 2206)) || ((pixel_index2 >= 2236) && (pixel_index2 <= 2238)) || ((pixel_index2 >= 2245) && (pixel_index2 <= 2246)) || pixel_index2 == 2250 || ((pixel_index2 >= 2252) && (pixel_index2 <= 2264)) || ((pixel_index2 >= 2274) && (pixel_index2 <= 2288)) || ((pixel_index2 >= 2291) && (pixel_index2 <= 2293)) || ((pixel_index2 >= 2296) && (pixel_index2 <= 2302)) || ((pixel_index2 >= 2332) && (pixel_index2 <= 2334)) || ((pixel_index2 >= 2341) && (pixel_index2 <= 2355)) || ((pixel_index2 >= 2374) && (pixel_index2 <= 2384)) || ((pixel_index2 >= 2392) && (pixel_index2 <= 2398)) || ((pixel_index2 >= 2428) && (pixel_index2 <= 2437)) || ((pixel_index2 >= 2443) && (pixel_index2 <= 2451)) || ((pixel_index2 >= 2470) && (pixel_index2 <= 2480)) || ((pixel_index2 >= 2487) && (pixel_index2 <= 2494)) || ((pixel_index2 >= 2526) && (pixel_index2 <= 2532)) || ((pixel_index2 >= 2540) && (pixel_index2 <= 2547)) || pixel_index2 == 2566 || ((pixel_index2 >= 2580) && (pixel_index2 <= 2588)) || ((pixel_index2 >= 2622) && (pixel_index2 <= 2626)) || pixel_index2 == 2636 || ((pixel_index2 >= 2639) && (pixel_index2 <= 2644)) || ((pixel_index2 >= 2647) && (pixel_index2 <= 2648)) || pixel_index2 == 2659 || ((pixel_index2 >= 2661) && (pixel_index2 <= 2662)) || ((pixel_index2 >= 2676) && (pixel_index2 <= 2684)) || ((pixel_index2 >= 2718) && (pixel_index2 <= 2721)) || pixel_index2 == 2732 || ((pixel_index2 >= 2735) && (pixel_index2 <= 2742)) || ((pixel_index2 >= 2756) && (pixel_index2 <= 2758)) || ((pixel_index2 >= 2772) && (pixel_index2 <= 2780)) || ((pixel_index2 >= 2814) && (pixel_index2 <= 2817)) || pixel_index2 == 2828 || ((pixel_index2 >= 2831) && (pixel_index2 <= 2838)) || ((pixel_index2 >= 2842) && (pixel_index2 <= 2848)) || ((pixel_index2 >= 2852) && (pixel_index2 <= 2859)) || ((pixel_index2 >= 2866) && (pixel_index2 <= 2876)) || ((pixel_index2 >= 2910) && (pixel_index2 <= 2913)) || pixel_index2 == 2924 || ((pixel_index2 >= 2927) && (pixel_index2 <= 2935)) || ((pixel_index2 >= 2938) && (pixel_index2 <= 2944)) || ((pixel_index2 >= 2947) && (pixel_index2 <= 2955)) || pixel_index2 == 2962 || ((pixel_index2 >= 2964) && (pixel_index2 <= 2972)) || ((pixel_index2 >= 3006) && (pixel_index2 <= 3013)) || ((pixel_index2 >= 3019) && (pixel_index2 <= 3021)) || ((pixel_index2 >= 3023) && (pixel_index2 <= 3032)) || ((pixel_index2 >= 3042) && (pixel_index2 <= 3051)) || ((pixel_index2 >= 3058) && (pixel_index2 <= 3060)) || pixel_index2 == 3063 || ((pixel_index2 >= 3065) && (pixel_index2 <= 3068)) || ((pixel_index2 >= 3102) && (pixel_index2 <= 3104)) || pixel_index2 == 3107 || ((pixel_index2 >= 3117) && (pixel_index2 <= 3123)) || ((pixel_index2 >= 3143) && (pixel_index2 <= 3147)) || ((pixel_index2 >= 3154) && (pixel_index2 <= 3155)) || pixel_index2 == 3159 || ((pixel_index2 >= 3161) && (pixel_index2 <= 3164)) || ((pixel_index2 >= 3198) && (pixel_index2 <= 3200)) || ((pixel_index2 >= 3202) && (pixel_index2 <= 3203)) || ((pixel_index2 >= 3213) && (pixel_index2 <= 3216)) || ((pixel_index2 >= 3218) && (pixel_index2 <= 3219)) || ((pixel_index2 >= 3239) && (pixel_index2 <= 3243)) || ((pixel_index2 >= 3250) && (pixel_index2 <= 3251)) || ((pixel_index2 >= 3255) && (pixel_index2 <= 3260)) || ((pixel_index2 >= 3292) && (pixel_index2 <= 3299)) || ((pixel_index2 >= 3309) && (pixel_index2 <= 3312)) || ((pixel_index2 >= 3314) && (pixel_index2 <= 3315)) || ((pixel_index2 >= 3335) && (pixel_index2 <= 3337)) || pixel_index2 == 3339 || ((pixel_index2 >= 3346) && (pixel_index2 <= 3347)) || ((pixel_index2 >= 3351) && (pixel_index2 <= 3352)) || ((pixel_index2 >= 3354) && (pixel_index2 <= 3358)) || ((pixel_index2 >= 3388) && (pixel_index2 <= 3393)) || pixel_index2 == 3395 || ((pixel_index2 >= 3405) && (pixel_index2 <= 3407)) || ((pixel_index2 >= 3409) && (pixel_index2 <= 3411)) || ((pixel_index2 >= 3431) && (pixel_index2 <= 3432)) || ((pixel_index2 >= 3434) && (pixel_index2 <= 3435)) || ((pixel_index2 >= 3438) && (pixel_index2 <= 3443)) || ((pixel_index2 >= 3447) && (pixel_index2 <= 3448)) || ((pixel_index2 >= 3450) && (pixel_index2 <= 3454)) || ((pixel_index2 >= 3484) && (pixel_index2 <= 3487)) || pixel_index2 == 3489 || pixel_index2 == 3491 || ((pixel_index2 >= 3501) && (pixel_index2 <= 3502)) || ((pixel_index2 >= 3505) && (pixel_index2 <= 3507)) || ((pixel_index2 >= 3527) && (pixel_index2 <= 3531)) || ((pixel_index2 >= 3538) && (pixel_index2 <= 3539)) || ((pixel_index2 >= 3543) && (pixel_index2 <= 3544)) || ((pixel_index2 >= 3546) && (pixel_index2 <= 3550)) || ((pixel_index2 >= 3580) && (pixel_index2 <= 3587)) || ((pixel_index2 >= 3597) && (pixel_index2 <= 3603)) || ((pixel_index2 >= 3623) && (pixel_index2 <= 3628)) || ((pixel_index2 >= 3633) && (pixel_index2 <= 3635)) || ((pixel_index2 >= 3639) && (pixel_index2 <= 3646)) || ((pixel_index2 >= 4620) && (pixel_index2 <= 4692)) || ((pixel_index2 >= 4707) && (pixel_index2 <= 4796)) || ((pixel_index2 >= 4803) && (pixel_index2 <= 4812)) || ((pixel_index2 >= 4814) && (pixel_index2 <= 4817)) || ((pixel_index2 >= 4819) && (pixel_index2 <= 4820)) || ((pixel_index2 >= 4827) && (pixel_index2 <= 4829)) || ((pixel_index2 >= 4834) && (pixel_index2 <= 4835)) || ((pixel_index2 >= 4838) && (pixel_index2 <= 4839)) || ((pixel_index2 >= 4841) && (pixel_index2 <= 4843)) || ((pixel_index2 >= 4845) && (pixel_index2 <= 4846)) || ((pixel_index2 >= 4851) && (pixel_index2 <= 4861)) || ((pixel_index2 >= 4863) && (pixel_index2 <= 4865)) || ((pixel_index2 >= 4868) && (pixel_index2 <= 4869)) || ((pixel_index2 >= 4871) && (pixel_index2 <= 4873)) || ((pixel_index2 >= 4880) && (pixel_index2 <= 4882)) || ((pixel_index2 >= 4887) && (pixel_index2 <= 4892)) || ((pixel_index2 >= 4899) && (pixel_index2 <= 4907)) || ((pixel_index2 >= 4910) && (pixel_index2 <= 4912)) || pixel_index2 == 4915 || pixel_index2 == 4924 || pixel_index2 == 4931 || pixel_index2 == 4935 || pixel_index2 == 4938 || pixel_index2 == 4941 || ((pixel_index2 >= 4948) && (pixel_index2 <= 4956)) || ((pixel_index2 >= 4959) && (pixel_index2 <= 4961)) || pixel_index2 == 4965 || pixel_index2 == 4968 || pixel_index2 == 4977 || ((pixel_index2 >= 4984) && (pixel_index2 <= 4988)) || ((pixel_index2 >= 4994) && (pixel_index2 <= 5003)) || ((pixel_index2 >= 5006) && (pixel_index2 <= 5008)) || pixel_index2 == 5011 || pixel_index2 == 5020 || pixel_index2 == 5027 || pixel_index2 == 5034 || pixel_index2 == 5037 || ((pixel_index2 >= 5044) && (pixel_index2 <= 5052)) || ((pixel_index2 >= 5055) && (pixel_index2 <= 5057)) || pixel_index2 == 5064 || pixel_index2 == 5073 || ((pixel_index2 >= 5080) && (pixel_index2 <= 5085)) || ((pixel_index2 >= 5090) && (pixel_index2 <= 5099)) || ((pixel_index2 >= 5102) && (pixel_index2 <= 5104)) || pixel_index2 == 5107 || ((pixel_index2 >= 5111) && (pixel_index2 <= 5112)) || ((pixel_index2 >= 5116) && (pixel_index2 <= 5119)) || ((pixel_index2 >= 5123) && (pixel_index2 <= 5124)) || pixel_index2 == 5130 || ((pixel_index2 >= 5133) && (pixel_index2 <= 5136)) || ((pixel_index2 >= 5140) && (pixel_index2 <= 5148)) || ((pixel_index2 >= 5151) && (pixel_index2 <= 5154)) || pixel_index2 == 5160 || ((pixel_index2 >= 5164) && (pixel_index2 <= 5165)) || pixel_index2 == 5169 || ((pixel_index2 >= 5173) && (pixel_index2 <= 5181)) || ((pixel_index2 >= 5186) && (pixel_index2 <= 5195)) || ((pixel_index2 >= 5198) && (pixel_index2 <= 5200)) || pixel_index2 == 5203 || ((pixel_index2 >= 5206) && (pixel_index2 <= 5209)) || ((pixel_index2 >= 5212) && (pixel_index2 <= 5216)) || ((pixel_index2 >= 5219) && (pixel_index2 <= 5220)) || pixel_index2 == 5226 || ((pixel_index2 >= 5229) && (pixel_index2 <= 5233)) || ((pixel_index2 >= 5236) && (pixel_index2 <= 5244)) || ((pixel_index2 >= 5247) && (pixel_index2 <= 5250)) || pixel_index2 == 5256 || ((pixel_index2 >= 5259) && (pixel_index2 <= 5262)) || pixel_index2 == 5265 || ((pixel_index2 >= 5271) && (pixel_index2 <= 5277)) || ((pixel_index2 >= 5282) && (pixel_index2 <= 5291)) || ((pixel_index2 >= 5294) && (pixel_index2 <= 5296)) || pixel_index2 == 5299 || ((pixel_index2 >= 5302) && (pixel_index2 <= 5305)) || ((pixel_index2 >= 5308) && (pixel_index2 <= 5312)) || pixel_index2 == 5315 || pixel_index2 == 5322 || ((pixel_index2 >= 5325) && (pixel_index2 <= 5329)) || ((pixel_index2 >= 5332) && (pixel_index2 <= 5340)) || ((pixel_index2 >= 5343) && (pixel_index2 <= 5345)) || pixel_index2 == 5352 || ((pixel_index2 >= 5355) && (pixel_index2 <= 5358)) || pixel_index2 == 5361 || ((pixel_index2 >= 5368) && (pixel_index2 <= 5373)) || ((pixel_index2 >= 5378) && (pixel_index2 <= 5387)) || ((pixel_index2 >= 5390) && (pixel_index2 <= 5392)) || pixel_index2 == 5395 || ((pixel_index2 >= 5398) && (pixel_index2 <= 5401)) || ((pixel_index2 >= 5404) && (pixel_index2 <= 5408)) || pixel_index2 == 5411 || pixel_index2 == 5415 || pixel_index2 == 5418 || ((pixel_index2 >= 5421) && (pixel_index2 <= 5425)) || ((pixel_index2 >= 5428) && (pixel_index2 <= 5436)) || ((pixel_index2 >= 5439) && (pixel_index2 <= 5441)) || pixel_index2 == 5445 || pixel_index2 == 5448 || ((pixel_index2 >= 5451) && (pixel_index2 <= 5454)) || ((pixel_index2 >= 5457) && (pixel_index2 <= 5458)) || ((pixel_index2 >= 5464) && (pixel_index2 <= 5469)) || ((pixel_index2 >= 5474) && (pixel_index2 <= 5483)) || ((pixel_index2 >= 5486) && (pixel_index2 <= 5488)) || pixel_index2 == 5491 || ((pixel_index2 >= 5494) && (pixel_index2 <= 5497)) || ((pixel_index2 >= 5500) && (pixel_index2 <= 5503)) || pixel_index2 == 5507 || ((pixel_index2 >= 5510) && (pixel_index2 <= 5511)) || pixel_index2 == 5514 || ((pixel_index2 >= 5517) && (pixel_index2 <= 5520)) || ((pixel_index2 >= 5524) && (pixel_index2 <= 5532)) || ((pixel_index2 >= 5535) && (pixel_index2 <= 5537)) || ((pixel_index2 >= 5540) && (pixel_index2 <= 5541)) || pixel_index2 == 5544 || ((pixel_index2 >= 5548) && (pixel_index2 <= 5549)) || ((pixel_index2 >= 5553) && (pixel_index2 <= 5556)) || ((pixel_index2 >= 5560) && (pixel_index2 <= 5565)) || ((pixel_index2 >= 5570) && (pixel_index2 <= 5575)) || pixel_index2 == 5584 || pixel_index2 == 5587 || ((pixel_index2 >= 5590) && (pixel_index2 <= 5593)) || pixel_index2 == 5596 || pixel_index2 == 5603 || pixel_index2 == 5610 || pixel_index2 == 5613 || ((pixel_index2 >= 5620) && (pixel_index2 <= 5624)) || pixel_index2 == 5633 || pixel_index2 == 5640 || pixel_index2 == 5649 || ((pixel_index2 >= 5656) && (pixel_index2 <= 5661)) || ((pixel_index2 >= 5667) && (pixel_index2 <= 5671)) || pixel_index2 == 5680 || pixel_index2 == 5683 || ((pixel_index2 >= 5686) && (pixel_index2 <= 5689)) || pixel_index2 == 5692 || pixel_index2 == 5699 || pixel_index2 == 5706 || pixel_index2 == 5709 || ((pixel_index2 >= 5716) && (pixel_index2 <= 5720)) || pixel_index2 == 5729 || pixel_index2 == 5736 || pixel_index2 == 5745 || ((pixel_index2 >= 5752) && (pixel_index2 <= 5756)) || ((pixel_index2 >= 5763) && (pixel_index2 <= 5768)) || ((pixel_index2 >= 5775) && (pixel_index2 <= 5776)) || ((pixel_index2 >= 5778) && (pixel_index2 <= 5780)) || ((pixel_index2 >= 5782) && (pixel_index2 <= 5785)) || ((pixel_index2 >= 5787) && (pixel_index2 <= 5789)) || ((pixel_index2 >= 5794) && (pixel_index2 <= 5796)) || ((pixel_index2 >= 5801) && (pixel_index2 <= 5802)) || ((pixel_index2 >= 5804) && (pixel_index2 <= 5806)) || ((pixel_index2 >= 5811) && (pixel_index2 <= 5817)) || ((pixel_index2 >= 5824) && (pixel_index2 <= 5826)) || ((pixel_index2 >= 5831) && (pixel_index2 <= 5833)) || ((pixel_index2 >= 5840) && (pixel_index2 <= 5842)) || ((pixel_index2 >= 5847) && (pixel_index2 <= 5852)) || (pixel_index2 >= 5868) && (pixel_index2 <= 5940)) oled_data2 = 16'b0000000000001010;
                    else if (pixel_index2 == 323 || pixel_index2 == 327 || pixel_index2 == 331 || pixel_index2 == 335 || pixel_index2 == 355 || pixel_index2 == 419 || pixel_index2 == 423 || pixel_index2 == 427 || pixel_index2 == 431 || pixel_index2 == 451 || pixel_index2 == 3253 || pixel_index2 == 3349) oled_data2 = 16'b0000010100000000;
                    else if (pixel_index2 == 511 || pixel_index2 == 531 || pixel_index2 == 535 || pixel_index2 == 539 || pixel_index2 == 543 || pixel_index2 == 551 || pixel_index2 == 555 || pixel_index2 == 559 || pixel_index2 == 563 || pixel_index2 == 567 || pixel_index2 == 571 || pixel_index2 == 607 || pixel_index2 == 627 || pixel_index2 == 631 || pixel_index2 == 635 || pixel_index2 == 639 || pixel_index2 == 647 || pixel_index2 == 651 || pixel_index2 == 655 || pixel_index2 == 659 || pixel_index2 == 663 || pixel_index2 == 667 || pixel_index2 == 3488) oled_data2 = 16'b1010000000000000;
                    else if (((pixel_index2 >= 895) && (pixel_index2 <= 896)) || ((pixel_index2 >= 899) && (pixel_index2 <= 900)) || ((pixel_index2 >= 903) && (pixel_index2 <= 904)) || ((pixel_index2 >= 907) && (pixel_index2 <= 908)) || ((pixel_index2 >= 911) && (pixel_index2 <= 912)) || ((pixel_index2 >= 915) && (pixel_index2 <= 916)) || ((pixel_index2 >= 919) && (pixel_index2 <= 920)) || ((pixel_index2 >= 923) && (pixel_index2 <= 924)) || ((pixel_index2 >= 927) && (pixel_index2 <= 928)) || ((pixel_index2 >= 931) && (pixel_index2 <= 932)) || ((pixel_index2 >= 935) && (pixel_index2 <= 936)) || ((pixel_index2 >= 939) && (pixel_index2 <= 940)) || ((pixel_index2 >= 943) && (pixel_index2 <= 944)) || ((pixel_index2 >= 947) && (pixel_index2 <= 948)) || ((pixel_index2 >= 951) && (pixel_index2 <= 952)) || ((pixel_index2 >= 955) && (pixel_index2 <= 956)) || pixel_index2 == 1155 || ((pixel_index2 >= 1159) && (pixel_index2 <= 1161)) || pixel_index2 == 1163 || ((pixel_index2 >= 1165) && (pixel_index2 <= 1166)) || pixel_index2 == 1168 || ((pixel_index2 >= 1170) && (pixel_index2 <= 1171)) || pixel_index2 == 1173 || ((pixel_index2 >= 1175) && (pixel_index2 <= 1176)) || pixel_index2 == 1254 || ((pixel_index2 >= 1256) && (pixel_index2 <= 1257)) || pixel_index2 == 1259 || ((pixel_index2 >= 1261) && (pixel_index2 <= 1262)) || ((pixel_index2 >= 1264) && (pixel_index2 <= 1267)) || ((pixel_index2 >= 1270) && (pixel_index2 <= 1272)) || pixel_index2 == 1350 || ((pixel_index2 >= 1352) && (pixel_index2 <= 1353)) || pixel_index2 == 1355 || ((pixel_index2 >= 1357) && (pixel_index2 <= 1358)) || pixel_index2 == 1360 || ((pixel_index2 >= 1362) && (pixel_index2 <= 1363)) || pixel_index2 == 1365 || ((pixel_index2 >= 1367) && (pixel_index2 <= 1368)) || ((pixel_index2 >= 1447) && (pixel_index2 <= 1449)) || ((pixel_index2 >= 1451) && (pixel_index2 <= 1454)) || ((pixel_index2 >= 1456) && (pixel_index2 <= 1459)) || ((pixel_index2 >= 1461) && (pixel_index2 <= 1464)) || pixel_index2 == 2213 || pixel_index2 == 2216 || ((pixel_index2 >= 2219) && (pixel_index2 <= 2221)) || pixel_index2 == 2223 || pixel_index2 == 2226 || ((pixel_index2 >= 2228) && (pixel_index2 <= 2230)) || pixel_index2 == 2310 || pixel_index2 == 2312 || pixel_index2 == 2314 || pixel_index2 == 2319 || pixel_index2 == 2322 || pixel_index2 == 2325 || ((pixel_index2 >= 2406) && (pixel_index2 <= 2408)) || ((pixel_index2 >= 2411) && (pixel_index2 <= 2412)) || ((pixel_index2 >= 2415) && (pixel_index2 <= 2416)) || pixel_index2 == 2418 || pixel_index2 == 2421 || pixel_index2 == 2501 || pixel_index2 == 2504 || pixel_index2 == 2509 || pixel_index2 == 2511 || ((pixel_index2 >= 2513) && (pixel_index2 <= 2514)) || pixel_index2 == 2517 || ((pixel_index2 >= 2598) && (pixel_index2 <= 2600)) || ((pixel_index2 >= 2602) && (pixel_index2 <= 2604)) || pixel_index2 == 2607 || pixel_index2 == 2610 || ((pixel_index2 >= 2612) && (pixel_index2 <= 2614)) || pixel_index2 == 2788 || pixel_index2 == 2791 || ((pixel_index2 >= 2794) && (pixel_index2 <= 2795)) || ((pixel_index2 >= 2799) && (pixel_index2 <= 2800)) || ((pixel_index2 >= 2804) && (pixel_index2 <= 2805)) || pixel_index2 == 2885 || pixel_index2 == 2887 || pixel_index2 == 2889 || pixel_index2 == 2892 || pixel_index2 == 2894 || pixel_index2 == 2897 || pixel_index2 == 2899 || pixel_index2 == 2902 || ((pixel_index2 >= 2982) && (pixel_index2 <= 2983)) || pixel_index2 == 2988 || pixel_index2 == 2990 || pixel_index2 == 2993 || pixel_index2 == 2998 || pixel_index2 == 3077 || pixel_index2 == 3079 || pixel_index2 == 3081 || pixel_index2 == 3084 || pixel_index2 == 3086 || pixel_index2 == 3089 || pixel_index2 == 3091 || pixel_index2 == 3094 || ((pixel_index2 >= 3133) && (pixel_index2 <= 3134)) || pixel_index2 == 3172 || pixel_index2 == 3175 || ((pixel_index2 >= 3178) && (pixel_index2 <= 3179)) || ((pixel_index2 >= 3183) && (pixel_index2 <= 3184)) || ((pixel_index2 >= 3188) && (pixel_index2 <= 3189)) || pixel_index2 == 3228 || pixel_index2 == 3327 || ((pixel_index2 >= 3364) && (pixel_index2 <= 3367)) || ((pixel_index2 >= 3370) && (pixel_index2 <= 3372)) || ((pixel_index2 >= 3375) && (pixel_index2 <= 3376)) || ((pixel_index2 >= 3380) && (pixel_index2 <= 3382)) || pixel_index2 == 3463 || pixel_index2 == 3465 || pixel_index2 == 3468 || pixel_index2 == 3470 || pixel_index2 == 3473 || pixel_index2 == 3475 || pixel_index2 == 3478 || pixel_index2 == 3559 || ((pixel_index2 >= 3562) && (pixel_index2 <= 3564)) || pixel_index2 == 3566 || pixel_index2 == 3569 || ((pixel_index2 >= 3572) && (pixel_index2 <= 3574)) || ((pixel_index2 >= 3630) && (pixel_index2 <= 3631)) || pixel_index2 == 3655 || pixel_index2 == 3657 || pixel_index2 == 3660 || pixel_index2 == 3662 || pixel_index2 == 3665 || pixel_index2 == 3667 || pixel_index2 == 3670 || pixel_index2 == 3751 || ((pixel_index2 >= 3754) && (pixel_index2 <= 3756)) || pixel_index2 == 3758 || pixel_index2 == 3761 || ((pixel_index2 >= 3764) && (pixel_index2 <= 3766)) || ((pixel_index2 >= 3938) && (pixel_index2 <= 3939)) || pixel_index2 == 3942 || pixel_index2 == 3945 || ((pixel_index2 >= 3947) && (pixel_index2 <= 3950)) || pixel_index2 == 3952 || ((pixel_index2 >= 3954) && (pixel_index2 <= 3955)) || ((pixel_index2 >= 3959) && (pixel_index2 <= 3962)) || ((pixel_index2 >= 3964) && (pixel_index2 <= 3967)) || ((pixel_index2 >= 3969) && (pixel_index2 <= 3972)) || ((pixel_index2 >= 3974) && (pixel_index2 <= 3977)) || pixel_index2 == 3979 || ((pixel_index2 >= 3981) && (pixel_index2 <= 3982)) || ((pixel_index2 >= 3984) && (pixel_index2 <= 3986)) || ((pixel_index2 >= 4008) && (pixel_index2 <= 4009)) || ((pixel_index2 >= 4012) && (pixel_index2 <= 4015)) || ((pixel_index2 >= 4017) && (pixel_index2 <= 4020)) || ((pixel_index2 >= 4022) && (pixel_index2 <= 4025)) || pixel_index2 == 4027 || ((pixel_index2 >= 4029) && (pixel_index2 <= 4030)) || ((pixel_index2 >= 4034) && (pixel_index2 <= 4035)) || ((pixel_index2 >= 4039) && (pixel_index2 <= 4040)) || ((pixel_index2 >= 4045) && (pixel_index2 <= 4046)) || pixel_index2 == 4048 || ((pixel_index2 >= 4050) && (pixel_index2 <= 4051)) || ((pixel_index2 >= 4057) && (pixel_index2 <= 4058)) || ((pixel_index2 >= 4060) && (pixel_index2 <= 4061)) || pixel_index2 == 4065 || ((pixel_index2 >= 4067) && (pixel_index2 <= 4068)) || pixel_index2 == 4070 || ((pixel_index2 >= 4072) && (pixel_index2 <= 4073)) || ((pixel_index2 >= 4075) && (pixel_index2 <= 4078)) || ((pixel_index2 >= 4082) && (pixel_index2 <= 4083)) || ((pixel_index2 >= 4104) && (pixel_index2 <= 4105)) || ((pixel_index2 >= 4110) && (pixel_index2 <= 4111)) || ((pixel_index2 >= 4113) && (pixel_index2 <= 4114)) || ((pixel_index2 >= 4120) && (pixel_index2 <= 4121)) || ((pixel_index2 >= 4124) && (pixel_index2 <= 4126)) || ((pixel_index2 >= 4130) && (pixel_index2 <= 4131)) || ((pixel_index2 >= 4135) && (pixel_index2 <= 4136)) || ((pixel_index2 >= 4139) && (pixel_index2 <= 4140)) || pixel_index2 == 4142 || pixel_index2 == 4144 || ((pixel_index2 >= 4146) && (pixel_index2 <= 4147)) || ((pixel_index2 >= 4151) && (pixel_index2 <= 4152)) || pixel_index2 == 4154 || ((pixel_index2 >= 4157) && (pixel_index2 <= 4159)) || pixel_index2 == 4161 || ((pixel_index2 >= 4163) && (pixel_index2 <= 4164)) || pixel_index2 == 4166 || ((pixel_index2 >= 4168) && (pixel_index2 <= 4169)) || pixel_index2 == 4171 || ((pixel_index2 >= 4173) && (pixel_index2 <= 4174)) || ((pixel_index2 >= 4178) && (pixel_index2 <= 4179)) || ((pixel_index2 >= 4200) && (pixel_index2 <= 4201)) || ((pixel_index2 >= 4204) && (pixel_index2 <= 4205)) || pixel_index2 == 4207 || ((pixel_index2 >= 4210) && (pixel_index2 <= 4212)) || ((pixel_index2 >= 4214) && (pixel_index2 <= 4215)) || pixel_index2 == 4217 || pixel_index2 == 4219 || ((pixel_index2 >= 4221) && (pixel_index2 <= 4222)) || ((pixel_index2 >= 4225) && (pixel_index2 <= 4228)) || pixel_index2 == 4230 || pixel_index2 == 4233 || ((pixel_index2 >= 4235) && (pixel_index2 <= 4238)) || ((pixel_index2 >= 4240) && (pixel_index2 <= 4243)) || ((pixel_index2 >= 4247) && (pixel_index2 <= 4250)) || ((pixel_index2 >= 4252) && (pixel_index2 <= 4254)) || ((pixel_index2 >= 4257) && (pixel_index2 <= 4260)) || ((pixel_index2 >= 4262) && (pixel_index2 <= 4265)) || pixel_index2 == 4267 || ((pixel_index2 >= 4269) && (pixel_index2 <= 4270)) || ((pixel_index2 >= 4272) && (pixel_index2 <= 4274)) || ((pixel_index2 >= 4295) && (pixel_index2 <= 4298)) || ((pixel_index2 >= 4300) && (pixel_index2 <= 4303)) || ((pixel_index2 >= 4305) && (pixel_index2 <= 4307)) || ((pixel_index2 >= 4310) && (pixel_index2 <= 4313)) || ((pixel_index2 >= 4315) && (pixel_index2 <= 4318)) || pixel_index2 == 4802 || pixel_index2 == 4893 || pixel_index2 == 5762 || pixel_index2 == 5853) oled_data2 = 16'b1111011110011110;
                    else if (pixel_index2 == 1086 || pixel_index2 == 1106 || pixel_index2 == 1110 || pixel_index2 == 1114 || pixel_index2 == 1118 || pixel_index2 == 1126 || pixel_index2 == 1130 || pixel_index2 == 1134 || pixel_index2 == 1138 || pixel_index2 == 1142 || pixel_index2 == 1146) oled_data2 = 16'b0000001010000000;
                    else if (pixel_index2 == 1090 || pixel_index2 == 1094 || pixel_index2 == 1098 || pixel_index2 == 1102 || pixel_index2 == 1122) oled_data2 = 16'b1111011110001010;
                    else if (((pixel_index2 >= 1190) && (pixel_index2 <= 1194)) || pixel_index2 == 1286 || pixel_index2 == 1290 || pixel_index2 == 1382 || pixel_index2 == 1386 || pixel_index2 == 1478 || pixel_index2 == 1482 || ((pixel_index2 >= 1574) && (pixel_index2 <= 1578)) || ((pixel_index2 >= 1637) && (pixel_index2 <= 1638)) || ((pixel_index2 >= 1641) && (pixel_index2 <= 1644)) || ((pixel_index2 >= 1646) && (pixel_index2 <= 1649)) || ((pixel_index2 >= 1652) && (pixel_index2 <= 1654)) || pixel_index2 == 1732 || pixel_index2 == 1735 || pixel_index2 == 1740 || pixel_index2 == 1745 || pixel_index2 == 1747 || pixel_index2 == 1753 || pixel_index2 == 1831 || pixel_index2 == 1836 || ((pixel_index2 >= 1839) && (pixel_index2 <= 1841)) || ((pixel_index2 >= 1844) && (pixel_index2 <= 1845)) || pixel_index2 == 1848 || pixel_index2 == 1924 || pixel_index2 == 1927 || pixel_index2 == 1932 || pixel_index2 == 1937 || pixel_index2 == 1942 || pixel_index2 == 1945 || ((pixel_index2 >= 2021) && (pixel_index2 <= 2022)) || pixel_index2 == 2028 || ((pixel_index2 >= 2030) && (pixel_index2 <= 2033)) || (pixel_index2 >= 2035) && (pixel_index2 <= 2037)) oled_data2 = 16'b0101010100011110;
                    else if (((pixel_index2 >= 1281) && (pixel_index2 <= 1282)) || pixel_index2 == 1292 || pixel_index2 == 1295 || ((pixel_index2 >= 1297) && (pixel_index2 <= 1299)) || pixel_index2 == 1302 || ((pixel_index2 >= 1304) && (pixel_index2 <= 1305)) || pixel_index2 == 1307 || pixel_index2 == 1309 || pixel_index2 == 1311 || pixel_index2 == 1313 || pixel_index2 == 1377 || ((pixel_index2 >= 1392) && (pixel_index2 <= 1395)) || ((pixel_index2 >= 1397) && (pixel_index2 <= 1399)) || pixel_index2 == 1401 || ((pixel_index2 >= 1403) && (pixel_index2 <= 1404)) || pixel_index2 == 1406 || pixel_index2 == 1409 || ((pixel_index2 >= 1487) && (pixel_index2 <= 1488)) || pixel_index2 == 1490 || pixel_index2 == 1493 || pixel_index2 == 1495 || pixel_index2 == 1497 || ((pixel_index2 >= 1499) && (pixel_index2 <= 1500)) || ((pixel_index2 >= 1502) && (pixel_index2 <= 1503)) || pixel_index2 == 1505 || pixel_index2 == 1697 || pixel_index2 == 1776 || ((pixel_index2 >= 1790) && (pixel_index2 <= 1791)) || pixel_index2 == 1793 || pixel_index2 == 1817 || pixel_index2 == 1871 || pixel_index2 == 1914 || pixel_index2 == 1974 || ((pixel_index2 >= 1989) && (pixel_index2 <= 1990)) || pixel_index2 == 1992 || pixel_index2 == 1995 || ((pixel_index2 >= 1997) && (pixel_index2 <= 1999)) || ((pixel_index2 >= 2009) && (pixel_index2 <= 2010)) || pixel_index2 == 2047 || ((pixel_index2 >= 2070) && (pixel_index2 <= 2071)) || pixel_index2 == 2083 || ((pixel_index2 >= 2086) && (pixel_index2 <= 2088)) || pixel_index2 == 2090 || pixel_index2 == 2094 || pixel_index2 == 2106 || pixel_index2 == 2141 || pixel_index2 == 2143 || ((pixel_index2 >= 2155) && (pixel_index2 <= 2156)) || pixel_index2 == 2179 || ((pixel_index2 >= 2185) && (pixel_index2 <= 2187)) || pixel_index2 == 2189 || pixel_index2 == 2240 || pixel_index2 == 2243 || pixel_index2 == 2251 || pixel_index2 == 2336 || pixel_index2 == 2338 || pixel_index2 == 2340 || pixel_index2 == 2548 || ((pixel_index2 >= 2550) && (pixel_index2 <= 2551)) || ((pixel_index2 >= 2562) && (pixel_index2 <= 2563)) || ((pixel_index2 >= 2567) && (pixel_index2 <= 2579)) || ((pixel_index2 >= 2645) && (pixel_index2 <= 2646)) || pixel_index2 == 2658 || pixel_index2 == 2660 || ((pixel_index2 >= 2663) && (pixel_index2 <= 2675)) || ((pixel_index2 >= 2759) && (pixel_index2 <= 2771)) || ((pixel_index2 >= 2925) && (pixel_index2 <= 2926)) || pixel_index2 == 2937 || pixel_index2 == 2946 || pixel_index2 == 3022 || ((pixel_index2 >= 3105) && (pixel_index2 <= 3106)) || pixel_index2 == 3201 || pixel_index2 == 3217 || ((pixel_index2 >= 3230) && (pixel_index2 <= 3231)) || pixel_index2 == 3313 || pixel_index2 == 3324 || pixel_index2 == 3408 || ((pixel_index2 >= 3421) && (pixel_index2 <= 3422)) || ((pixel_index2 >= 3503) && (pixel_index2 <= 3504)) || ((pixel_index2 >= 3533) && (pixel_index2 <= 3536)) || pixel_index2 == 3629 || pixel_index2 == 3632) oled_data2 = 16'b1010010100010100;
                    else if (pixel_index2 == 1287 || pixel_index2 == 1289 || pixel_index2 == 1479 || pixel_index2 == 1481 || pixel_index2 == 1667 || pixel_index2 == 1669 || pixel_index2 == 1671 || pixel_index2 == 1673 || pixel_index2 == 1675 || pixel_index2 == 1677 || pixel_index2 == 1859 || pixel_index2 == 1861 || pixel_index2 == 1863 || pixel_index2 == 1865 || pixel_index2 == 1867 || pixel_index2 == 1869 || ((pixel_index2 >= 1879) && (pixel_index2 <= 1881)) || ((pixel_index2 >= 1889) && (pixel_index2 <= 1891)) || ((pixel_index2 >= 1975) && (pixel_index2 <= 1987)) || ((pixel_index2 >= 2002) && (pixel_index2 <= 2007)) || pixel_index2 == 2055 || pixel_index2 == 2057 || ((pixel_index2 >= 2072) && (pixel_index2 <= 2073)) || ((pixel_index2 >= 2081) && (pixel_index2 <= 2082)) || ((pixel_index2 >= 2097) && (pixel_index2 <= 2103)) || pixel_index2 == 2169 || pixel_index2 == 2177 || ((pixel_index2 >= 2193) && (pixel_index2 <= 2194)) || ((pixel_index2 >= 2198) && (pixel_index2 <= 2199)) || pixel_index2 == 2239 || ((pixel_index2 >= 2241) && (pixel_index2 <= 2242)) || pixel_index2 == 2244 || pixel_index2 == 2247 || pixel_index2 == 2249 || pixel_index2 == 2265 || pixel_index2 == 2273 || ((pixel_index2 >= 2289) && (pixel_index2 <= 2290)) || ((pixel_index2 >= 2294) && (pixel_index2 <= 2295)) || pixel_index2 == 2335 || pixel_index2 == 2337 || pixel_index2 == 2339 || ((pixel_index2 >= 2356) && (pixel_index2 <= 2361)) || ((pixel_index2 >= 2369) && (pixel_index2 <= 2373)) || ((pixel_index2 >= 2385) && (pixel_index2 <= 2391)) || ((pixel_index2 >= 2438) && (pixel_index2 <= 2442)) || ((pixel_index2 >= 2452) && (pixel_index2 <= 2457)) || ((pixel_index2 >= 2465) && (pixel_index2 <= 2469)) || ((pixel_index2 >= 2481) && (pixel_index2 <= 2486)) || pixel_index2 == 2533 || pixel_index2 == 2539 || pixel_index2 == 2549 || ((pixel_index2 >= 2552) && (pixel_index2 <= 2553)) || pixel_index2 == 2561 || ((pixel_index2 >= 2564) && (pixel_index2 <= 2565)) || ((pixel_index2 >= 2627) && (pixel_index2 <= 2629)) || pixel_index2 == 2635 || ((pixel_index2 >= 2637) && (pixel_index2 <= 2638)) || pixel_index2 == 2649 || pixel_index2 == 2657 || ((pixel_index2 >= 2722) && (pixel_index2 <= 2725)) || pixel_index2 == 2731 || ((pixel_index2 >= 2733) && (pixel_index2 <= 2734)) || ((pixel_index2 >= 2743) && (pixel_index2 <= 2755)) || ((pixel_index2 >= 2818) && (pixel_index2 <= 2821)) || pixel_index2 == 2827 || ((pixel_index2 >= 2829) && (pixel_index2 <= 2830)) || ((pixel_index2 >= 2839) && (pixel_index2 <= 2841)) || ((pixel_index2 >= 2849) && (pixel_index2 <= 2851)) || ((pixel_index2 >= 2914) && (pixel_index2 <= 2917)) || pixel_index2 == 2923 || pixel_index2 == 2936 || pixel_index2 == 2945 || pixel_index2 == 2963 || ((pixel_index2 >= 3014) && (pixel_index2 <= 3018)) || ((pixel_index2 >= 3061) && (pixel_index2 <= 3062)) || pixel_index2 == 3064 || ((pixel_index2 >= 3108) && (pixel_index2 <= 3116)) || pixel_index2 == 3160 || ((pixel_index2 >= 3204) && (pixel_index2 <= 3212)) || ((pixel_index2 >= 3300) && (pixel_index2 <= 3308)) || pixel_index2 == 3317 || ((pixel_index2 >= 3319) && (pixel_index2 <= 3320)) || ((pixel_index2 >= 3330) && (pixel_index2 <= 3331)) || pixel_index2 == 3333 || pixel_index2 == 3338 || ((pixel_index2 >= 3396) && (pixel_index2 <= 3404)) || pixel_index2 == 3433 || ((pixel_index2 >= 3436) && (pixel_index2 <= 3437)) || ((pixel_index2 >= 3492) && (pixel_index2 <= 3500)) || ((pixel_index2 >= 3588) && (pixel_index2 <= 3596)) || ((pixel_index2 >= 3684) && (pixel_index2 <= 3692)) || ((pixel_index2 >= 3724) && (pixel_index2 <= 3729)) || ((pixel_index2 >= 3820) && (pixel_index2 <= 3825)) || ((pixel_index2 >= 3893) && (pixel_index2 <= 3894)) || ((pixel_index2 >= 3897) && (pixel_index2 <= 3905)) || ((pixel_index2 >= 3908) && (pixel_index2 <= 3909)) || ((pixel_index2 >= 3989) && (pixel_index2 <= 3990)) || ((pixel_index2 >= 3994) && (pixel_index2 <= 4000)) || ((pixel_index2 >= 4004) && (pixel_index2 <= 4005)) || ((pixel_index2 >= 4085) && (pixel_index2 <= 4086)) || ((pixel_index2 >= 4090) && (pixel_index2 <= 4096)) || ((pixel_index2 >= 4100) && (pixel_index2 <= 4101)) || pixel_index2 == 4706 || pixel_index2 == 4797 || pixel_index2 == 5666 || pixel_index2 == 5757) oled_data2 = 16'b0101001010001010;
                    else if (pixel_index2 == 1296 || ((pixel_index2 >= 1300) && (pixel_index2 <= 1301)) || pixel_index2 == 1303 || pixel_index2 == 1306 || pixel_index2 == 1308 || pixel_index2 == 1310 || pixel_index2 == 1312 || pixel_index2 == 1391 || pixel_index2 == 1396 || pixel_index2 == 1400 || pixel_index2 == 1402 || pixel_index2 == 1405 || ((pixel_index2 >= 1407) && (pixel_index2 <= 1408)) || pixel_index2 == 1489 || ((pixel_index2 >= 1491) && (pixel_index2 <= 1492)) || pixel_index2 == 1494 || pixel_index2 == 1496 || pixel_index2 == 1498 || pixel_index2 == 1501 || pixel_index2 == 1504 || pixel_index2 == 3353 || pixel_index2 == 3449 || pixel_index2 == 3545) oled_data2 = 16'b0101001010010100;
                    else if (((pixel_index2 >= 1317) && (pixel_index2 <= 1319)) || ((pixel_index2 >= 1322) && (pixel_index2 <= 1324)) || ((pixel_index2 >= 1327) && (pixel_index2 <= 1329)) || ((pixel_index2 >= 1332) && (pixel_index2 <= 1334)) || pixel_index2 == 1415 || pixel_index2 == 1420 || pixel_index2 == 1425 || pixel_index2 == 1428 || pixel_index2 == 1511 || pixel_index2 == 1516 || ((pixel_index2 >= 1519) && (pixel_index2 <= 1521)) || ((pixel_index2 >= 1524) && (pixel_index2 <= 1526)) || pixel_index2 == 1607 || pixel_index2 == 1612 || pixel_index2 == 1617 || pixel_index2 == 1622 || ((pixel_index2 >= 1701) && (pixel_index2 <= 1703)) || pixel_index2 == 1708 || ((pixel_index2 >= 1711) && (pixel_index2 <= 1713)) || (pixel_index2 >= 1716) && (pixel_index2 <= 1718)) oled_data2 = 16'b1010000000001010;
                    else if (pixel_index2 == 3229 || (pixel_index2 >= 3325) && (pixel_index2 <= 3326)) oled_data2 = 16'b0101010100001010;
                    else if (pixel_index2 == 3394 || pixel_index2 == 3490) oled_data2 = 16'b0000000000010100;
                    else if (pixel_index2 == 3532 || pixel_index2 == 3537) oled_data2 = 16'b0101000000000000;
                    else if (((pixel_index2 >= 4423) && (pixel_index2 <= 4505)) || ((pixel_index2 >= 4513) && (pixel_index2 <= 4518)) || (pixel_index2 >= 4602) && (pixel_index2 <= 4606)) oled_data2 = 16'b0000001010011110;
                    else if (((pixel_index2 >= 4519) && (pixel_index2 <= 4601)) || ((pixel_index2 >= 4609) && (pixel_index2 <= 4619)) || ((pixel_index2 >= 4693) && (pixel_index2 <= 4702)) || pixel_index2 == 4705 || pixel_index2 == 4798 || pixel_index2 == 4801 || pixel_index2 == 4894 || ((pixel_index2 >= 4897) && (pixel_index2 <= 4898)) || ((pixel_index2 >= 4989) && (pixel_index2 <= 4990)) || pixel_index2 == 4993 || pixel_index2 == 5086 || pixel_index2 == 5089 || pixel_index2 == 5182 || pixel_index2 == 5185 || pixel_index2 == 5278 || pixel_index2 == 5281 || pixel_index2 == 5374 || pixel_index2 == 5377 || pixel_index2 == 5470 || pixel_index2 == 5473 || pixel_index2 == 5566 || pixel_index2 == 5569 || pixel_index2 == 5662 || pixel_index2 == 5665 || pixel_index2 == 5758 || pixel_index2 == 5761 || pixel_index2 == 5854 || ((pixel_index2 >= 5857) && (pixel_index2 <= 5867)) || ((pixel_index2 >= 5941) && (pixel_index2 <= 5950)) || (pixel_index2 >= 5959) && (pixel_index2 <= 6041)) oled_data2 = 16'b0000001010010100;
                    else if (pixel_index2 == 4813 || pixel_index2 == 4818 || ((pixel_index2 >= 4821) && (pixel_index2 <= 4826)) || ((pixel_index2 >= 4830) && (pixel_index2 <= 4833)) || ((pixel_index2 >= 4836) && (pixel_index2 <= 4837)) || pixel_index2 == 4840 || pixel_index2 == 4844 || ((pixel_index2 >= 4847) && (pixel_index2 <= 4850)) || pixel_index2 == 4862 || ((pixel_index2 >= 4866) && (pixel_index2 <= 4867)) || pixel_index2 == 4870 || ((pixel_index2 >= 4874) && (pixel_index2 <= 4879)) || ((pixel_index2 >= 4883) && (pixel_index2 <= 4886)) || pixel_index2 == 4908 || pixel_index2 == 4913 || pixel_index2 == 4916 || pixel_index2 == 4923 || pixel_index2 == 4925 || pixel_index2 == 4930 || pixel_index2 == 4934 || pixel_index2 == 4937 || pixel_index2 == 4939 || pixel_index2 == 4942 || pixel_index2 == 4947 || pixel_index2 == 4957 || pixel_index2 == 4964 || pixel_index2 == 4967 || pixel_index2 == 4969 || pixel_index2 == 4976 || pixel_index2 == 4978 || pixel_index2 == 4983 || pixel_index2 == 5031 || pixel_index2 == 5061 || pixel_index2 == 5221 || pixel_index2 == 5251 || ((pixel_index2 >= 5268) && (pixel_index2 <= 5270)) || pixel_index2 == 5316 || pixel_index2 == 5346 || pixel_index2 == 5367 || pixel_index2 == 5504 || pixel_index2 == 5521 || pixel_index2 == 5547 || pixel_index2 == 5550 || pixel_index2 == 5557 || ((pixel_index2 >= 5576) && (pixel_index2 <= 5579)) || ((pixel_index2 >= 5582) && (pixel_index2 <= 5583)) || ((pixel_index2 >= 5597) && (pixel_index2 <= 5599)) || ((pixel_index2 >= 5606) && (pixel_index2 <= 5607)) || ((pixel_index2 >= 5614) && (pixel_index2 <= 5616)) || ((pixel_index2 >= 5625) && (pixel_index2 <= 5628)) || ((pixel_index2 >= 5631) && (pixel_index2 <= 5632)) || ((pixel_index2 >= 5636) && (pixel_index2 <= 5637)) || ((pixel_index2 >= 5644) && (pixel_index2 <= 5645)) || (pixel_index2 >= 5650) && (pixel_index2 <= 5652)) oled_data2 = 16'b0101001010000000;
                    else if (pixel_index2 == 4909 || pixel_index2 == 4914 || ((pixel_index2 >= 4917) && (pixel_index2 <= 4922)) || ((pixel_index2 >= 4926) && (pixel_index2 <= 4929)) || ((pixel_index2 >= 4932) && (pixel_index2 <= 4933)) || pixel_index2 == 4936 || pixel_index2 == 4940 || ((pixel_index2 >= 4943) && (pixel_index2 <= 4946)) || pixel_index2 == 4958 || ((pixel_index2 >= 4962) && (pixel_index2 <= 4963)) || pixel_index2 == 4966 || ((pixel_index2 >= 4970) && (pixel_index2 <= 4975)) || ((pixel_index2 >= 4979) && (pixel_index2 <= 4982)) || ((pixel_index2 >= 5004) && (pixel_index2 <= 5005)) || ((pixel_index2 >= 5009) && (pixel_index2 <= 5010)) || ((pixel_index2 >= 5012) && (pixel_index2 <= 5019)) || ((pixel_index2 >= 5021) && (pixel_index2 <= 5026)) || ((pixel_index2 >= 5028) && (pixel_index2 <= 5030)) || ((pixel_index2 >= 5032) && (pixel_index2 <= 5033)) || ((pixel_index2 >= 5035) && (pixel_index2 <= 5036)) || ((pixel_index2 >= 5038) && (pixel_index2 <= 5043)) || ((pixel_index2 >= 5053) && (pixel_index2 <= 5054)) || ((pixel_index2 >= 5058) && (pixel_index2 <= 5060)) || ((pixel_index2 >= 5062) && (pixel_index2 <= 5063)) || ((pixel_index2 >= 5065) && (pixel_index2 <= 5072)) || ((pixel_index2 >= 5074) && (pixel_index2 <= 5079)) || ((pixel_index2 >= 5100) && (pixel_index2 <= 5101)) || ((pixel_index2 >= 5105) && (pixel_index2 <= 5106)) || ((pixel_index2 >= 5108) && (pixel_index2 <= 5110)) || ((pixel_index2 >= 5113) && (pixel_index2 <= 5115)) || ((pixel_index2 >= 5120) && (pixel_index2 <= 5122)) || ((pixel_index2 >= 5125) && (pixel_index2 <= 5129)) || ((pixel_index2 >= 5131) && (pixel_index2 <= 5132)) || ((pixel_index2 >= 5137) && (pixel_index2 <= 5139)) || ((pixel_index2 >= 5149) && (pixel_index2 <= 5150)) || ((pixel_index2 >= 5155) && (pixel_index2 <= 5159)) || ((pixel_index2 >= 5161) && (pixel_index2 <= 5163)) || ((pixel_index2 >= 5166) && (pixel_index2 <= 5168)) || ((pixel_index2 >= 5170) && (pixel_index2 <= 5172)) || ((pixel_index2 >= 5196) && (pixel_index2 <= 5197)) || ((pixel_index2 >= 5201) && (pixel_index2 <= 5202)) || ((pixel_index2 >= 5204) && (pixel_index2 <= 5205)) || ((pixel_index2 >= 5210) && (pixel_index2 <= 5211)) || ((pixel_index2 >= 5217) && (pixel_index2 <= 5218)) || ((pixel_index2 >= 5222) && (pixel_index2 <= 5225)) || ((pixel_index2 >= 5227) && (pixel_index2 <= 5228)) || ((pixel_index2 >= 5234) && (pixel_index2 <= 5235)) || ((pixel_index2 >= 5245) && (pixel_index2 <= 5246)) || ((pixel_index2 >= 5252) && (pixel_index2 <= 5255)) || ((pixel_index2 >= 5257) && (pixel_index2 <= 5258)) || ((pixel_index2 >= 5263) && (pixel_index2 <= 5264)) || ((pixel_index2 >= 5266) && (pixel_index2 <= 5267)) || ((pixel_index2 >= 5292) && (pixel_index2 <= 5293)) || ((pixel_index2 >= 5297) && (pixel_index2 <= 5298)) || ((pixel_index2 >= 5300) && (pixel_index2 <= 5301)) || ((pixel_index2 >= 5306) && (pixel_index2 <= 5307)) || ((pixel_index2 >= 5313) && (pixel_index2 <= 5314)) || ((pixel_index2 >= 5317) && (pixel_index2 <= 5321)) || ((pixel_index2 >= 5323) && (pixel_index2 <= 5324)) || ((pixel_index2 >= 5330) && (pixel_index2 <= 5331)) || ((pixel_index2 >= 5341) && (pixel_index2 <= 5342)) || ((pixel_index2 >= 5347) && (pixel_index2 <= 5351)) || ((pixel_index2 >= 5353) && (pixel_index2 <= 5354)) || ((pixel_index2 >= 5359) && (pixel_index2 <= 5360)) || ((pixel_index2 >= 5362) && (pixel_index2 <= 5366)) || ((pixel_index2 >= 5388) && (pixel_index2 <= 5389)) || ((pixel_index2 >= 5393) && (pixel_index2 <= 5394)) || ((pixel_index2 >= 5396) && (pixel_index2 <= 5397)) || ((pixel_index2 >= 5402) && (pixel_index2 <= 5403)) || ((pixel_index2 >= 5409) && (pixel_index2 <= 5410)) || ((pixel_index2 >= 5412) && (pixel_index2 <= 5414)) || ((pixel_index2 >= 5416) && (pixel_index2 <= 5417)) || ((pixel_index2 >= 5419) && (pixel_index2 <= 5420)) || ((pixel_index2 >= 5426) && (pixel_index2 <= 5427)) || ((pixel_index2 >= 5437) && (pixel_index2 <= 5438)) || ((pixel_index2 >= 5442) && (pixel_index2 <= 5444)) || ((pixel_index2 >= 5446) && (pixel_index2 <= 5447)) || ((pixel_index2 >= 5449) && (pixel_index2 <= 5450)) || ((pixel_index2 >= 5455) && (pixel_index2 <= 5456)) || ((pixel_index2 >= 5459) && (pixel_index2 <= 5463)) || ((pixel_index2 >= 5484) && (pixel_index2 <= 5485)) || ((pixel_index2 >= 5489) && (pixel_index2 <= 5490)) || ((pixel_index2 >= 5492) && (pixel_index2 <= 5493)) || ((pixel_index2 >= 5498) && (pixel_index2 <= 5499)) || ((pixel_index2 >= 5505) && (pixel_index2 <= 5506)) || ((pixel_index2 >= 5508) && (pixel_index2 <= 5509)) || ((pixel_index2 >= 5512) && (pixel_index2 <= 5513)) || ((pixel_index2 >= 5515) && (pixel_index2 <= 5516)) || ((pixel_index2 >= 5522) && (pixel_index2 <= 5523)) || ((pixel_index2 >= 5533) && (pixel_index2 <= 5534)) || ((pixel_index2 >= 5538) && (pixel_index2 <= 5539)) || ((pixel_index2 >= 5542) && (pixel_index2 <= 5543)) || ((pixel_index2 >= 5545) && (pixel_index2 <= 5546)) || ((pixel_index2 >= 5551) && (pixel_index2 <= 5552)) || ((pixel_index2 >= 5558) && (pixel_index2 <= 5559)) || ((pixel_index2 >= 5580) && (pixel_index2 <= 5581)) || ((pixel_index2 >= 5585) && (pixel_index2 <= 5586)) || ((pixel_index2 >= 5588) && (pixel_index2 <= 5589)) || ((pixel_index2 >= 5594) && (pixel_index2 <= 5595)) || ((pixel_index2 >= 5600) && (pixel_index2 <= 5602)) || ((pixel_index2 >= 5604) && (pixel_index2 <= 5605)) || ((pixel_index2 >= 5608) && (pixel_index2 <= 5609)) || ((pixel_index2 >= 5611) && (pixel_index2 <= 5612)) || ((pixel_index2 >= 5617) && (pixel_index2 <= 5619)) || ((pixel_index2 >= 5629) && (pixel_index2 <= 5630)) || ((pixel_index2 >= 5634) && (pixel_index2 <= 5635)) || ((pixel_index2 >= 5638) && (pixel_index2 <= 5639)) || ((pixel_index2 >= 5641) && (pixel_index2 <= 5643)) || ((pixel_index2 >= 5646) && (pixel_index2 <= 5648)) || ((pixel_index2 >= 5653) && (pixel_index2 <= 5655)) || ((pixel_index2 >= 5672) && (pixel_index2 <= 5679)) || ((pixel_index2 >= 5681) && (pixel_index2 <= 5682)) || ((pixel_index2 >= 5684) && (pixel_index2 <= 5685)) || ((pixel_index2 >= 5690) && (pixel_index2 <= 5691)) || ((pixel_index2 >= 5693) && (pixel_index2 <= 5698)) || ((pixel_index2 >= 5700) && (pixel_index2 <= 5705)) || ((pixel_index2 >= 5707) && (pixel_index2 <= 5708)) || ((pixel_index2 >= 5710) && (pixel_index2 <= 5715)) || ((pixel_index2 >= 5721) && (pixel_index2 <= 5728)) || ((pixel_index2 >= 5730) && (pixel_index2 <= 5735)) || ((pixel_index2 >= 5737) && (pixel_index2 <= 5744)) || ((pixel_index2 >= 5746) && (pixel_index2 <= 5751)) || ((pixel_index2 >= 5769) && (pixel_index2 <= 5774)) || pixel_index2 == 5777 || pixel_index2 == 5781 || pixel_index2 == 5786 || ((pixel_index2 >= 5790) && (pixel_index2 <= 5793)) || ((pixel_index2 >= 5797) && (pixel_index2 <= 5800)) || pixel_index2 == 5803 || ((pixel_index2 >= 5807) && (pixel_index2 <= 5810)) || ((pixel_index2 >= 5818) && (pixel_index2 <= 5823)) || ((pixel_index2 >= 5827) && (pixel_index2 <= 5830)) || ((pixel_index2 >= 5834) && (pixel_index2 <= 5839)) || (pixel_index2 >= 5843) && (pixel_index2 <= 5846)) oled_data2 = 16'b1111010100010100;
                    else oled_data2 = 0;
                end
            endcase
           
    end
    if (sorting_algorithm == 4'b0001) begin // bubble sorting
        // 2nd OLED
        if (((pixel_index2 >= 0) && (pixel_index2 <= 96)) || ((pixel_index2 >= 191) && (pixel_index2 <= 192)) || ((pixel_index2 >= 287) && (pixel_index2 <= 288)) || ((pixel_index2 >= 383) && (pixel_index2 <= 384)) || ((pixel_index2 >= 479) && (pixel_index2 <= 480)) || ((pixel_index2 >= 575) && (pixel_index2 <= 576)) || ((pixel_index2 >= 671) && (pixel_index2 <= 672)) || ((pixel_index2 >= 767) && (pixel_index2 <= 768)) || ((pixel_index2 >= 863) && (pixel_index2 <= 864)) || ((pixel_index2 >= 959) && (pixel_index2 <= 960)) || ((pixel_index2 >= 1055) && (pixel_index2 <= 1056)) || ((pixel_index2 >= 1151) && (pixel_index2 <= 1152)) || ((pixel_index2 >= 1247) && (pixel_index2 <= 1248)) || ((pixel_index2 >= 1343) && (pixel_index2 <= 1344)) || ((pixel_index2 >= 1439) && (pixel_index2 <= 1440)) || ((pixel_index2 >= 1535) && (pixel_index2 <= 1536)) || ((pixel_index2 >= 1631) && (pixel_index2 <= 1632)) || ((pixel_index2 >= 1727) && (pixel_index2 <= 1728)) || ((pixel_index2 >= 1823) && (pixel_index2 <= 1824)) || ((pixel_index2 >= 1919) && (pixel_index2 <= 1920)) || ((pixel_index2 >= 2015) && (pixel_index2 <= 2016)) || ((pixel_index2 >= 2111) && (pixel_index2 <= 2112)) || ((pixel_index2 >= 2207) && (pixel_index2 <= 2208)) || ((pixel_index2 >= 2303) && (pixel_index2 <= 2304)) || ((pixel_index2 >= 2399) && (pixel_index2 <= 2400)) || ((pixel_index2 >= 2495) && (pixel_index2 <= 2496)) || ((pixel_index2 >= 2591) && (pixel_index2 <= 2592)) || ((pixel_index2 >= 2687) && (pixel_index2 <= 2688)) || ((pixel_index2 >= 2783) && (pixel_index2 <= 2784)) || ((pixel_index2 >= 2879) && (pixel_index2 <= 2880)) || ((pixel_index2 >= 2975) && (pixel_index2 <= 2976)) || ((pixel_index2 >= 3071) && (pixel_index2 <= 3072)) || ((pixel_index2 >= 3167) && (pixel_index2 <= 3168)) || ((pixel_index2 >= 3263) && (pixel_index2 <= 3264)) || ((pixel_index2 >= 3359) && (pixel_index2 <= 3360)) || ((pixel_index2 >= 3455) && (pixel_index2 <= 3456)) || ((pixel_index2 >= 3551) && (pixel_index2 <= 3552)) || ((pixel_index2 >= 3647) && (pixel_index2 <= 3743)) || ((pixel_index2 >= 4050) && (pixel_index2 <= 4054)) || ((pixel_index2 >= 4058) && (pixel_index2 <= 4062)) || ((pixel_index2 >= 4147) && (pixel_index2 <= 4150)) || ((pixel_index2 >= 4154) && (pixel_index2 <= 4158)) || pixel_index2 == 4242 || ((pixel_index2 >= 4245) && (pixel_index2 <= 4246)) || ((pixel_index2 >= 4250) && (pixel_index2 <= 4254)) || pixel_index2 == 4339 || ((pixel_index2 >= 4341) && (pixel_index2 <= 4342)) || ((pixel_index2 >= 4346) && (pixel_index2 <= 4349)) || pixel_index2 == 4434 || pixel_index2 == 4436 || pixel_index2 == 4438 || ((pixel_index2 >= 4442) && (pixel_index2 <= 4443)) || pixel_index2 == 4446 || pixel_index2 == 4530 || pixel_index2 == 4532 || pixel_index2 == 4534 || pixel_index2 == 4538 || ((pixel_index2 >= 4540) && (pixel_index2 <= 4542)) || ((pixel_index2 >= 4626) && (pixel_index2 <= 4628)) || pixel_index2 == 4630 || ((pixel_index2 >= 4635) && (pixel_index2 <= 4638)) || ((pixel_index2 >= 4722) && (pixel_index2 <= 4723)) || ((pixel_index2 >= 4725) && (pixel_index2 <= 4726)) || ((pixel_index2 >= 4730) && (pixel_index2 <= 4734)) || pixel_index2 == 4818 || ((pixel_index2 >= 4821) && (pixel_index2 <= 4822)) || ((pixel_index2 >= 4826) && (pixel_index2 <= 4830)) || ((pixel_index2 >= 4915) && (pixel_index2 <= 4918)) || ((pixel_index2 >= 4922) && (pixel_index2 <= 4926)) || ((pixel_index2 >= 5010) && (pixel_index2 <= 5014)) || ((pixel_index2 >= 5019) && (pixel_index2 <= 5022)) || ((pixel_index2 >= 5106) && (pixel_index2 <= 5110)) || ((pixel_index2 >= 5116) && (pixel_index2 <= 5118)) || ((pixel_index2 >= 5202) && (pixel_index2 <= 5206)) || ((pixel_index2 >= 5212) && (pixel_index2 <= 5214)) || ((pixel_index2 >= 5309) && (pixel_index2 <= 5310)) || pixel_index2 == 5402 || ((pixel_index2 >= 5405) && (pixel_index2 <= 5406)) || pixel_index2 == 5498 || pixel_index2 == 5595 || pixel_index2 == 5690 || (pixel_index2 >= 5692) && (pixel_index2 <= 5693)) oled_data2 = 16'b1111010100000000;
        else if (pixel_index2 == 440 || ((pixel_index2 >= 442) && (pixel_index2 <= 443)) || ((pixel_index2 >= 446) && (pixel_index2 <= 447)) || pixel_index2 == 450 || pixel_index2 == 455 || pixel_index2 == 458 || ((pixel_index2 >= 462) && (pixel_index2 <= 463)) || pixel_index2 == 469 || pixel_index2 == 471 || pixel_index2 == 473 || pixel_index2 == 475 || pixel_index2 == 538 || pixel_index2 == 540 || pixel_index2 == 544 || pixel_index2 == 547 || pixel_index2 == 551 || pixel_index2 == 553 || pixel_index2 == 555 || pixel_index2 == 557 || pixel_index2 == 565 || pixel_index2 == 567 || pixel_index2 == 569 || pixel_index2 == 572 || pixel_index2 == 634 || pixel_index2 == 636 || ((pixel_index2 >= 638) && (pixel_index2 <= 640)) || pixel_index2 == 643 || pixel_index2 == 645 || pixel_index2 == 647 || pixel_index2 == 649 || pixel_index2 == 651 || ((pixel_index2 >= 654) && (pixel_index2 <= 655)) || pixel_index2 == 661 || pixel_index2 == 663 || pixel_index2 == 665 || pixel_index2 == 668 || ((pixel_index2 >= 730) && (pixel_index2 <= 731)) || pixel_index2 == 735 || ((pixel_index2 >= 738) && (pixel_index2 <= 739)) || pixel_index2 == 742 || pixel_index2 == 746 || ((pixel_index2 >= 749) && (pixel_index2 <= 750)) || pixel_index2 == 757 || pixel_index2 == 759 || pixel_index2 == 761 || ((pixel_index2 >= 763) && (pixel_index2 <= 764)) || pixel_index2 == 826 || pixel_index2 == 835 || pixel_index2 == 853 || pixel_index2 == 855 || pixel_index2 == 860 || pixel_index2 == 922 || pixel_index2 == 931 || pixel_index2 == 949 || pixel_index2 == 951 || pixel_index2 == 953 || pixel_index2 == 956 || pixel_index2 == 1018 || pixel_index2 == 1027 || pixel_index2 == 1045 || pixel_index2 == 1047 || pixel_index2 == 1052 || pixel_index2 == 1387 || pixel_index2 == 1482 || pixel_index2 == 1484 || pixel_index2 == 1519 || pixel_index2 == 1578 || pixel_index2 == 1615 || ((pixel_index2 >= 1635) && (pixel_index2 <= 1636)) || pixel_index2 == 1638 || pixel_index2 == 1641 || pixel_index2 == 1643 || ((pixel_index2 >= 1645) && (pixel_index2 <= 1646)) || pixel_index2 == 1649 || pixel_index2 == 1653 || ((pixel_index2 >= 1655) && (pixel_index2 <= 1656)) || pixel_index2 == 1659 || ((pixel_index2 >= 1661) && (pixel_index2 <= 1662)) || ((pixel_index2 >= 1674) && (pixel_index2 <= 1675)) || ((pixel_index2 >= 1679) && (pixel_index2 <= 1680)) || pixel_index2 == 1684 || ((pixel_index2 >= 1686) && (pixel_index2 <= 1687)) || ((pixel_index2 >= 1690) && (pixel_index2 <= 1691)) || pixel_index2 == 1694 || pixel_index2 == 1696 || ((pixel_index2 >= 1706) && (pixel_index2 <= 1707)) || ((pixel_index2 >= 1710) && (pixel_index2 <= 1711)) || ((pixel_index2 >= 1713) && (pixel_index2 <= 1714)) || pixel_index2 == 1718 || pixel_index2 == 1720 || ((pixel_index2 >= 1724) && (pixel_index2 <= 1725)) || pixel_index2 == 1730 || pixel_index2 == 1735 || pixel_index2 == 1737 || pixel_index2 == 1739 || pixel_index2 == 1743 || pixel_index2 == 1745 || pixel_index2 == 1747 || pixel_index2 == 1749 || pixel_index2 == 1753 || pixel_index2 == 1755 || pixel_index2 == 1759 || pixel_index2 == 1770 || pixel_index2 == 1772 || pixel_index2 == 1774 || pixel_index2 == 1776 || pixel_index2 == 1780 || pixel_index2 == 1782 || pixel_index2 == 1784 || pixel_index2 == 1788 || pixel_index2 == 1790 || pixel_index2 == 1792 || pixel_index2 == 1801 || pixel_index2 == 1805 || pixel_index2 == 1807 || pixel_index2 == 1809 || pixel_index2 == 1811 || pixel_index2 == 1813 || pixel_index2 == 1815 || pixel_index2 == 1817 || pixel_index2 == 1819 || ((pixel_index2 >= 1827) && (pixel_index2 <= 1828)) || pixel_index2 == 1831 || pixel_index2 == 1833 || pixel_index2 == 1835 || ((pixel_index2 >= 1837) && (pixel_index2 <= 1839)) || pixel_index2 == 1841 || pixel_index2 == 1843 || pixel_index2 == 1845 || ((pixel_index2 >= 1847) && (pixel_index2 <= 1849)) || pixel_index2 == 1851 || ((pixel_index2 >= 1853) && (pixel_index2 <= 1855)) || pixel_index2 == 1866 || pixel_index2 == 1868 || pixel_index2 == 1870 || pixel_index2 == 1872 || pixel_index2 == 1874 || pixel_index2 == 1876 || pixel_index2 == 1878 || pixel_index2 == 1880 || ((pixel_index2 >= 1882) && (pixel_index2 <= 1884)) || pixel_index2 == 1886 || pixel_index2 == 1888 || ((pixel_index2 >= 1898) && (pixel_index2 <= 1899)) || pixel_index2 == 1901 || pixel_index2 == 1903 || pixel_index2 == 1905 || pixel_index2 == 1907 || pixel_index2 == 1909 || pixel_index2 == 1911 || pixel_index2 == 1913 || ((pixel_index2 >= 1916) && (pixel_index2 <= 1917)) || ((pixel_index2 >= 1922) && (pixel_index2 <= 1923)) || ((pixel_index2 >= 1926) && (pixel_index2 <= 1927)) || ((pixel_index2 >= 1930) && (pixel_index2 <= 1931)) || pixel_index2 == 1934 || pixel_index2 == 1938 || ((pixel_index2 >= 1940) && (pixel_index2 <= 1941)) || pixel_index2 == 1944 || pixel_index2 == 1947 || pixel_index2 == 1950 || pixel_index2 == 1962 || pixel_index2 == 1964 || ((pixel_index2 >= 1967) && (pixel_index2 <= 1968)) || ((pixel_index2 >= 1971) && (pixel_index2 <= 1972)) || pixel_index2 == 1975 || pixel_index2 == 1979 || ((pixel_index2 >= 1983) && (pixel_index2 <= 1984)) || ((pixel_index2 >= 1993) && (pixel_index2 <= 1994)) || ((pixel_index2 >= 1998) && (pixel_index2 <= 1999)) || pixel_index2 == 2002 || pixel_index2 == 2005 || pixel_index2 == 2009 || ((pixel_index2 >= 2011) && (pixel_index2 <= 2012)) || pixel_index2 == 2023 || pixel_index2 == 2043 || pixel_index2 == 2064 || pixel_index2 == 2119 || pixel_index2 == 2139 || pixel_index2 == 2160 || pixel_index2 == 2215 || pixel_index2 == 2235 || pixel_index2 == 2256 || pixel_index2 == 2645 || pixel_index2 == 2692 || pixel_index2 == 2740 || pixel_index2 == 2742 || pixel_index2 == 2787 || pixel_index2 == 2836 || pixel_index2 == 2883 || pixel_index2 == 2886 || pixel_index2 == 2888 || pixel_index2 == 2891 || pixel_index2 == 2894 || pixel_index2 == 2896 || ((pixel_index2 >= 2899) && (pixel_index2 <= 2900)) || ((pixel_index2 >= 2903) && (pixel_index2 <= 2904)) || pixel_index2 == 2909 || pixel_index2 == 2911 || ((pixel_index2 >= 2913) && (pixel_index2 <= 2914)) || ((pixel_index2 >= 2923) && (pixel_index2 <= 2925)) || ((pixel_index2 >= 2932) && (pixel_index2 <= 2933)) || pixel_index2 == 2936 || pixel_index2 == 2938 || pixel_index2 == 2940 || pixel_index2 == 2943 || ((pixel_index2 >= 2951) && (pixel_index2 <= 2952)) || ((pixel_index2 >= 2954) && (pixel_index2 <= 2955)) || ((pixel_index2 >= 2959) && (pixel_index2 <= 2960)) || ((pixel_index2 >= 2963) && (pixel_index2 <= 2964)) || ((pixel_index2 >= 2966) && (pixel_index2 <= 2967)) || pixel_index2 == 2973 || pixel_index2 == 2982 || pixel_index2 == 2984 || pixel_index2 == 2986 || pixel_index2 == 2988 || pixel_index2 == 2990 || pixel_index2 == 2993 || pixel_index2 == 2997 || pixel_index2 == 3001 || pixel_index2 == 3005 || pixel_index2 == 3007 || pixel_index2 == 3009 || pixel_index2 == 3011 || pixel_index2 == 3020 || pixel_index2 == 3028 || pixel_index2 == 3030 || pixel_index2 == 3032 || pixel_index2 == 3034 || pixel_index2 == 3036 || pixel_index2 == 3038 || pixel_index2 == 3040 || pixel_index2 == 3046 || pixel_index2 == 3052 || pixel_index2 == 3054 || pixel_index2 == 3058 || pixel_index2 == 3062 || pixel_index2 == 3064 || pixel_index2 == 3069 || pixel_index2 == 3078 || pixel_index2 == 3080 || pixel_index2 == 3082 || pixel_index2 == 3084 || pixel_index2 == 3086 || pixel_index2 == 3089 || pixel_index2 == 3093 || ((pixel_index2 >= 3095) && (pixel_index2 <= 3097)) || pixel_index2 == 3099 || pixel_index2 == 3101 || pixel_index2 == 3103 || pixel_index2 == 3105 || pixel_index2 == 3107 || pixel_index2 == 3116 || pixel_index2 == 3124 || pixel_index2 == 3126 || pixel_index2 == 3128 || pixel_index2 == 3130 || pixel_index2 == 3132 || pixel_index2 == 3134 || pixel_index2 == 3136 || ((pixel_index2 >= 3143) && (pixel_index2 <= 3144)) || ((pixel_index2 >= 3146) && (pixel_index2 <= 3148)) || ((pixel_index2 >= 3151) && (pixel_index2 <= 3152)) || ((pixel_index2 >= 3155) && (pixel_index2 <= 3156)) || pixel_index2 == 3158 || pixel_index2 == 3160 || pixel_index2 == 3165 || ((pixel_index2 >= 3175) && (pixel_index2 <= 3176)) || pixel_index2 == 3179 || pixel_index2 == 3182 || ((pixel_index2 >= 3184) && (pixel_index2 <= 3185)) || ((pixel_index2 >= 3187) && (pixel_index2 <= 3188)) || pixel_index2 == 3192 || ((pixel_index2 >= 3196) && (pixel_index2 <= 3197)) || pixel_index2 == 3199 || ((pixel_index2 >= 3201) && (pixel_index2 <= 3202)) || pixel_index2 == 3212 || pixel_index2 == 3220 || pixel_index2 == 3222 || pixel_index2 == 3224 || ((pixel_index2 >= 3227) && (pixel_index2 <= 3228)) || pixel_index2 == 3231 || ((pixel_index2 >= 3238) && (pixel_index2 <= 3239)) || pixel_index2 == 3243 || ((pixel_index2 >= 3246) && (pixel_index2 <= 3247)) || ((pixel_index2 >= 3250) && (pixel_index2 <= 3251)) || pixel_index2 == 3255 || ((pixel_index2 >= 3259) && (pixel_index2 <= 3261)) || pixel_index2 == 3281 || pixel_index2 == 3297 || pixel_index2 == 3308 || pixel_index2 == 3320 || pixel_index2 == 3354 || pixel_index2 == 3357 || pixel_index2 == 3374 || pixel_index2 == 3377 || pixel_index2 == 3391 || pixel_index2 == 3393 || ((pixel_index2 >= 3404) && (pixel_index2 <= 3405)) || pixel_index2 == 3416 || pixel_index2 == 3450 || pixel_index2 == 3453 || pixel_index2 == 3473 || pixel_index2 == 3489 || pixel_index2 == 3500 || pixel_index2 == 3512 || ((pixel_index2 >= 3547) && (pixel_index2 <= 3549)) || ((pixel_index2 >= 3840) && (pixel_index2 <= 3936)) || ((pixel_index2 >= 4031) && (pixel_index2 <= 4032)) || ((pixel_index2 >= 4103) && (pixel_index2 <= 4104)) || pixel_index2 == 4110 || ((pixel_index2 >= 4114) && (pixel_index2 <= 4116)) || ((pixel_index2 >= 4120) && (pixel_index2 <= 4123)) || ((pixel_index2 >= 4127) && (pixel_index2 <= 4128)) || pixel_index2 == 4198 || pixel_index2 == 4200 || pixel_index2 == 4206 || pixel_index2 == 4209 || pixel_index2 == 4213 || ((pixel_index2 >= 4215) && (pixel_index2 <= 4216)) || ((pixel_index2 >= 4219) && (pixel_index2 <= 4220)) || ((pixel_index2 >= 4223) && (pixel_index2 <= 4224)) || ((pixel_index2 >= 4243) && (pixel_index2 <= 4244)) || pixel_index2 == 4296 || pixel_index2 == 4302 || pixel_index2 == 4305 || pixel_index2 == 4309 || ((pixel_index2 >= 4311) && (pixel_index2 <= 4312)) || ((pixel_index2 >= 4319) && (pixel_index2 <= 4320)) || pixel_index2 == 4340 || ((pixel_index2 >= 4351) && (pixel_index2 <= 4352)) || pixel_index2 == 4354 || pixel_index2 == 4392 || pixel_index2 == 4395 || pixel_index2 == 4398 || pixel_index2 == 4401 || pixel_index2 == 4405 || ((pixel_index2 >= 4407) && (pixel_index2 <= 4408)) || ((pixel_index2 >= 4415) && (pixel_index2 <= 4416)) || pixel_index2 == 4437 || ((pixel_index2 >= 4451) && (pixel_index2 <= 4452)) || ((pixel_index2 >= 4486) && (pixel_index2 <= 4489)) || ((pixel_index2 >= 4492) && (pixel_index2 <= 4493)) || pixel_index2 == 4495 || ((pixel_index2 >= 4498) && (pixel_index2 <= 4500)) || ((pixel_index2 >= 4504) && (pixel_index2 <= 4506)) || ((pixel_index2 >= 4511) && (pixel_index2 <= 4512)) || pixel_index2 == 4525 || pixel_index2 == 4549 || pixel_index2 == 4584 || ((pixel_index2 >= 4602) && (pixel_index2 <= 4603)) || ((pixel_index2 >= 4607) && (pixel_index2 <= 4608)) || pixel_index2 == 4612 || pixel_index2 == 4621 || pixel_index2 == 4646 || pixel_index2 == 4680 || ((pixel_index2 >= 4699) && (pixel_index2 <= 4700)) || ((pixel_index2 >= 4703) && (pixel_index2 <= 4704)) || pixel_index2 == 4709 || pixel_index2 == 4718 || pixel_index2 == 4743 || pixel_index2 == 4776 || ((pixel_index2 >= 4791) && (pixel_index2 <= 4792)) || ((pixel_index2 >= 4795) && (pixel_index2 <= 4796)) || ((pixel_index2 >= 4799) && (pixel_index2 <= 4800)) || ((pixel_index2 >= 4814) && (pixel_index2 <= 4815)) || pixel_index2 == 4839 || pixel_index2 == 4872 || ((pixel_index2 >= 4888) && (pixel_index2 <= 4891)) || ((pixel_index2 >= 4895) && (pixel_index2 <= 4897)) || pixel_index2 == 4913 || pixel_index2 == 4936 || ((pixel_index2 >= 4991) && (pixel_index2 <= 4992)) || pixel_index2 == 4994 || pixel_index2 == 5016 || ((pixel_index2 >= 5087) && (pixel_index2 <= 5088)) || pixel_index2 == 5101 || pixel_index2 == 5112 || pixel_index2 == 5128 || ((pixel_index2 >= 5149) && (pixel_index2 <= 5152)) || pixel_index2 == 5155 || ((pixel_index2 >= 5158) && (pixel_index2 <= 5161)) || ((pixel_index2 >= 5164) && (pixel_index2 <= 5167)) || ((pixel_index2 >= 5169) && (pixel_index2 <= 5172)) || ((pixel_index2 >= 5176) && (pixel_index2 <= 5180)) || ((pixel_index2 >= 5183) && (pixel_index2 <= 5184)) || pixel_index2 == 5199 || pixel_index2 == 5224 || pixel_index2 == 5249 || pixel_index2 == 5251 || pixel_index2 == 5253 || pixel_index2 == 5257 || pixel_index2 == 5259 || pixel_index2 == 5263 || pixel_index2 == 5265 || pixel_index2 == 5269 || pixel_index2 == 5271 || pixel_index2 == 5276 || ((pixel_index2 >= 5279) && (pixel_index2 <= 5280)) || pixel_index2 == 5296 || pixel_index2 == 5304 || ((pixel_index2 >= 5341) && (pixel_index2 <= 5345)) || pixel_index2 == 5347 || pixel_index2 == 5349 || pixel_index2 == 5353 || pixel_index2 == 5355 || pixel_index2 == 5359 || pixel_index2 == 5361 || pixel_index2 == 5365 || pixel_index2 == 5367 || pixel_index2 == 5372 || ((pixel_index2 >= 5375) && (pixel_index2 <= 5376)) || pixel_index2 == 5401 || pixel_index2 == 5437 || pixel_index2 == 5441 || pixel_index2 == 5443 || pixel_index2 == 5445 || pixel_index2 == 5449 || pixel_index2 == 5451 || pixel_index2 == 5455 || pixel_index2 == 5457 || pixel_index2 == 5461 || pixel_index2 == 5463 || pixel_index2 == 5468 || ((pixel_index2 >= 5471) && (pixel_index2 <= 5472)) || pixel_index2 == 5489 || pixel_index2 == 5497 || ((pixel_index2 >= 5534) && (pixel_index2 <= 5536)) || pixel_index2 == 5539 || ((pixel_index2 >= 5542) && (pixel_index2 <= 5545)) || ((pixel_index2 >= 5548) && (pixel_index2 <= 5551)) || pixel_index2 == 5553 || pixel_index2 == 5557 || ((pixel_index2 >= 5560) && (pixel_index2 <= 5564)) || ((pixel_index2 >= 5567) && (pixel_index2 <= 5568)) || pixel_index2 == 5575 || pixel_index2 == 5585 || pixel_index2 == 5594 || pixel_index2 == 5635 || pixel_index2 == 5641 || pixel_index2 == 5647 || pixel_index2 == 5657 || pixel_index2 == 5660 || ((pixel_index2 >= 5663) && (pixel_index2 <= 5664)) || pixel_index2 == 5691 || pixel_index2 == 5731 || pixel_index2 == 5737 || pixel_index2 == 5743 || pixel_index2 == 5752 || pixel_index2 == 5756 || ((pixel_index2 >= 5759) && (pixel_index2 <= 5760)) || pixel_index2 == 5767 || pixel_index2 == 5789 || pixel_index2 == 5827 || pixel_index2 == 5833 || pixel_index2 == 5839 || pixel_index2 == 5848 || pixel_index2 == 5852 || ((pixel_index2 >= 5855) && (pixel_index2 <= 5856)) || pixel_index2 == 5864 || ((pixel_index2 >= 5886) && (pixel_index2 <= 5888)) || pixel_index2 == 5890 || pixel_index2 == 5923 || pixel_index2 == 5929 || pixel_index2 == 5935 || ((pixel_index2 >= 5945) && (pixel_index2 <= 5948)) || ((pixel_index2 >= 5951) && (pixel_index2 <= 5952)) || pixel_index2 == 5961 || ((pixel_index2 >= 6047) && (pixel_index2 <= 6059)) || pixel_index2 == 6061 || (pixel_index2 >= 6063) && (pixel_index2 <= 6143)) oled_data2 = 16'b1111011110011110;
        else if (((pixel_index2 >= 4042) && (pixel_index2 <= 4046)) || ((pixel_index2 >= 4138) && (pixel_index2 <= 4142)) || ((pixel_index2 >= 4234) && (pixel_index2 <= 4237)) || ((pixel_index2 >= 4330) && (pixel_index2 <= 4333)) || ((pixel_index2 >= 4426) && (pixel_index2 <= 4428)) || pixel_index2 == 4430 || ((pixel_index2 >= 4522) && (pixel_index2 <= 4524)) || pixel_index2 == 4526 || ((pixel_index2 >= 4618) && (pixel_index2 <= 4620)) || pixel_index2 == 4622 || ((pixel_index2 >= 4714) && (pixel_index2 <= 4717)) || ((pixel_index2 >= 4810) && (pixel_index2 <= 4813)) || (pixel_index2 >= 4906) && (pixel_index2 <= 4910)) oled_data2 = 16'b1010000000000000;
        else if (((pixel_index2 >= 4066) && (pixel_index2 <= 4070)) || ((pixel_index2 >= 4162) && (pixel_index2 <= 4166)) || ((pixel_index2 >= 4258) && (pixel_index2 <= 4262)) || ((pixel_index2 >= 4355) && (pixel_index2 <= 4358)) || pixel_index2 == 4450 || ((pixel_index2 >= 4453) && (pixel_index2 <= 4454)) || ((pixel_index2 >= 4547) && (pixel_index2 <= 4548)) || pixel_index2 == 4550 || pixel_index2 == 4645) oled_data2 = 16'b0000010100000000;
        else if (((pixel_index2 >= 4144) && (pixel_index2 <= 4146)) || ((pixel_index2 >= 4238) && (pixel_index2 <= 4239)) || pixel_index2 == 4334 || pixel_index2 == 4350 || pixel_index2 == 4353 || pixel_index2 == 4429 || ((pixel_index2 >= 4444) && (pixel_index2 <= 4445)) || pixel_index2 == 4533 || pixel_index2 == 4539 || ((pixel_index2 >= 4610) && (pixel_index2 <= 4611)) || pixel_index2 == 4629 || pixel_index2 == 4634 || pixel_index2 == 4705 || pixel_index2 == 4724 || pixel_index2 == 4729 || pixel_index2 == 4801 || pixel_index2 == 4805 || ((pixel_index2 >= 4819) && (pixel_index2 <= 4820)) || pixel_index2 == 4825 || pixel_index2 == 4901 || pixel_index2 == 4912 || pixel_index2 == 4914 || pixel_index2 == 4920 || ((pixel_index2 >= 4995) && (pixel_index2 <= 4996)) || pixel_index2 == 5032 || ((pixel_index2 >= 5098) && (pixel_index2 <= 5100)) || pixel_index2 == 5102 || pixel_index2 == 5193 || pixel_index2 == 5208 || pixel_index2 == 5288 || pixel_index2 == 5320 || pixel_index2 == 5383 || pixel_index2 == 5393 || pixel_index2 == 5415 || pixel_index2 == 5479 || pixel_index2 == 5511 || pixel_index2 == 5606 || pixel_index2 == 5671 || pixel_index2 == 5681 || pixel_index2 == 5701 || pixel_index2 == 5777 || pixel_index2 == 5788 || ((pixel_index2 >= 5795) && (pixel_index2 <= 5796)) || pixel_index2 == 5872 || pixel_index2 == 5889 || pixel_index2 == 5967 || pixel_index2 == 6060 || pixel_index2 == 6062) oled_data2 = 16'b0101001010001010;
        else if (((pixel_index2 >= 4337) && (pixel_index2 <= 4338)) || pixel_index2 == 4435 || pixel_index2 == 4527 || pixel_index2 == 4531 || ((pixel_index2 >= 4544) && (pixel_index2 <= 4545)) || pixel_index2 == 4624 || pixel_index2 == 4642 || pixel_index2 == 4708 || pixel_index2 == 4721 || pixel_index2 == 4933 || pixel_index2 == 5018 || pixel_index2 == 5030 || pixel_index2 == 5114 || pixel_index2 == 5126 || pixel_index2 == 5210 || pixel_index2 == 5293 || pixel_index2 == 5307 || pixel_index2 == 5487 || pixel_index2 == 5598 || pixel_index2 == 5673 || ((pixel_index2 >= 5695) && (pixel_index2 <= 5697)) || pixel_index2 == 5867) oled_data2 = 16'b0101010100011110;
        else if (pixel_index2 == 4543 || pixel_index2 == 4739 || pixel_index2 == 4836 || pixel_index2 == 5115 || pixel_index2 == 5211 || pixel_index2 == 5222 || pixel_index2 == 5308 || pixel_index2 == 5502 || pixel_index2 == 5577 || ((pixel_index2 >= 5599) && (pixel_index2 <= 5600)) || pixel_index2 == 5868) oled_data2 = 16'b1010001010011110;
        else if (pixel_index2 == 4546 || pixel_index2 == 4623 || ((pixel_index2 >= 4643) && (pixel_index2 <= 4644)) || pixel_index2 == 4720 || pixel_index2 == 4741 || pixel_index2 == 4837 || pixel_index2 == 4898 || pixel_index2 == 4934 || pixel_index2 == 5294 || pixel_index2 == 5306 || pixel_index2 == 5391 || pixel_index2 == 5403 || ((pixel_index2 >= 5499) && (pixel_index2 <= 5500)) || ((pixel_index2 >= 5596) && (pixel_index2 <= 5597)) || pixel_index2 == 5694 || pixel_index2 == 5769 || pixel_index2 == 5866) oled_data2 = 16'b1010010100011110;
        else if (pixel_index2 == 4740 || pixel_index2 == 5390 || pixel_index2 == 5770) oled_data2 = 16'b0101000000010100;
        else if (pixel_index2 == 5404 || pixel_index2 == 5501) oled_data2 = 16'b1010000000011110;
        else oled_data2 = 0;
    end 
    else if (sorting_algorithm == 4'b0010) begin // selection sorting
        if (((pixel_index2 >= 0) && (pixel_index2 <= 96)) || ((pixel_index2 >= 191) && (pixel_index2 <= 192)) || ((pixel_index2 >= 287) && (pixel_index2 <= 288)) || ((pixel_index2 >= 383) && (pixel_index2 <= 384)) || ((pixel_index2 >= 479) && (pixel_index2 <= 480)) || ((pixel_index2 >= 575) && (pixel_index2 <= 576)) || ((pixel_index2 >= 671) && (pixel_index2 <= 672)) || ((pixel_index2 >= 767) && (pixel_index2 <= 768)) || ((pixel_index2 >= 863) && (pixel_index2 <= 864)) || ((pixel_index2 >= 959) && (pixel_index2 <= 960)) || ((pixel_index2 >= 1055) && (pixel_index2 <= 1056)) || ((pixel_index2 >= 1151) && (pixel_index2 <= 1152)) || ((pixel_index2 >= 1247) && (pixel_index2 <= 1248)) || ((pixel_index2 >= 1343) && (pixel_index2 <= 1344)) || ((pixel_index2 >= 1439) && (pixel_index2 <= 1440)) || ((pixel_index2 >= 1535) && (pixel_index2 <= 1536)) || ((pixel_index2 >= 1631) && (pixel_index2 <= 1632)) || ((pixel_index2 >= 1727) && (pixel_index2 <= 1728)) || ((pixel_index2 >= 1823) && (pixel_index2 <= 1824)) || ((pixel_index2 >= 1919) && (pixel_index2 <= 1920)) || ((pixel_index2 >= 2015) && (pixel_index2 <= 2016)) || ((pixel_index2 >= 2111) && (pixel_index2 <= 2112)) || ((pixel_index2 >= 2207) && (pixel_index2 <= 2208)) || ((pixel_index2 >= 2303) && (pixel_index2 <= 2304)) || ((pixel_index2 >= 2399) && (pixel_index2 <= 2400)) || ((pixel_index2 >= 2495) && (pixel_index2 <= 2496)) || ((pixel_index2 >= 2591) && (pixel_index2 <= 2592)) || ((pixel_index2 >= 2687) && (pixel_index2 <= 2688)) || ((pixel_index2 >= 2783) && (pixel_index2 <= 2784)) || ((pixel_index2 >= 2879) && (pixel_index2 <= 2880)) || ((pixel_index2 >= 2975) && (pixel_index2 <= 2976)) || ((pixel_index2 >= 3071) && (pixel_index2 <= 3072)) || ((pixel_index2 >= 3167) && (pixel_index2 <= 3168)) || ((pixel_index2 >= 3263) && (pixel_index2 <= 3264)) || ((pixel_index2 >= 3359) && (pixel_index2 <= 3360)) || ((pixel_index2 >= 3455) && (pixel_index2 <= 3456)) || ((pixel_index2 >= 3551) && (pixel_index2 <= 3552)) || ((pixel_index2 >= 3647) && (pixel_index2 <= 3743)) || ((pixel_index2 >= 4145) && (pixel_index2 <= 4149)) || ((pixel_index2 >= 4241) && (pixel_index2 <= 4245)) || ((pixel_index2 >= 4337) && (pixel_index2 <= 4341)) || ((pixel_index2 >= 4433) && (pixel_index2 <= 4437)) || ((pixel_index2 >= 4529) && (pixel_index2 <= 4533)) || ((pixel_index2 >= 4625) && (pixel_index2 <= 4629)) || ((pixel_index2 >= 4722) && (pixel_index2 <= 4725)) || ((pixel_index2 >= 4818) && (pixel_index2 <= 4821)) || ((pixel_index2 >= 4914) && (pixel_index2 <= 4917)) || ((pixel_index2 >= 5011) && (pixel_index2 <= 5013)) || ((pixel_index2 >= 5107) && (pixel_index2 <= 5109)) || ((pixel_index2 >= 5203) && (pixel_index2 <= 5205)) || ((pixel_index2 >= 5300) && (pixel_index2 <= 5301)) || ((pixel_index2 >= 5396) && (pixel_index2 <= 5397)) || ((pixel_index2 >= 5492) && (pixel_index2 <= 5493)) || pixel_index2 == 5585 || ((pixel_index2 >= 5588) && (pixel_index2 <= 5589)) || ((pixel_index2 >= 5681) && (pixel_index2 <= 5685)) || (pixel_index2 >= 5777) && (pixel_index2 <= 5781)) oled_data2 = 16'b1111010100000000;
        else if (pixel_index2 == 249 || pixel_index2 == 345 || pixel_index2 == 386 || ((pixel_index2 >= 388) && (pixel_index2 <= 389)) || ((pixel_index2 >= 392) && (pixel_index2 <= 393)) || pixel_index2 == 396 || pixel_index2 == 401 || pixel_index2 == 404 || ((pixel_index2 >= 408) && (pixel_index2 <= 409)) || pixel_index2 == 415 || pixel_index2 == 417 || pixel_index2 == 419 || pixel_index2 == 421 || pixel_index2 == 428 || ((pixel_index2 >= 431) && (pixel_index2 <= 432)) || ((pixel_index2 >= 435) && (pixel_index2 <= 436)) || ((pixel_index2 >= 440) && (pixel_index2 <= 441)) || ((pixel_index2 >= 443) && (pixel_index2 <= 444)) || pixel_index2 == 447 || pixel_index2 == 451 || pixel_index2 == 459 || pixel_index2 == 461 || pixel_index2 == 464 || pixel_index2 == 466 || pixel_index2 == 469 || pixel_index2 == 474 || pixel_index2 == 477 || pixel_index2 == 484 || pixel_index2 == 486 || pixel_index2 == 490 || pixel_index2 == 493 || pixel_index2 == 497 || pixel_index2 == 499 || pixel_index2 == 501 || pixel_index2 == 503 || pixel_index2 == 511 || pixel_index2 == 513 || pixel_index2 == 515 || pixel_index2 == 518 || pixel_index2 == 525 || pixel_index2 == 527 || pixel_index2 == 529 || pixel_index2 == 533 || pixel_index2 == 535 || pixel_index2 == 537 || pixel_index2 == 541 || pixel_index2 == 543 || pixel_index2 == 547 || pixel_index2 == 558 || pixel_index2 == 560 || pixel_index2 == 562 || pixel_index2 == 564 || pixel_index2 == 566 || pixel_index2 == 570 || pixel_index2 == 573 || pixel_index2 == 580 || pixel_index2 == 582 || ((pixel_index2 >= 584) && (pixel_index2 <= 586)) || pixel_index2 == 589 || pixel_index2 == 591 || pixel_index2 == 593 || pixel_index2 == 595 || pixel_index2 == 597 || ((pixel_index2 >= 600) && (pixel_index2 <= 601)) || pixel_index2 == 607 || pixel_index2 == 609 || pixel_index2 == 611 || pixel_index2 == 614 || pixel_index2 == 621 || pixel_index2 == 623 || pixel_index2 == 625 || ((pixel_index2 >= 627) && (pixel_index2 <= 629)) || pixel_index2 == 631 || pixel_index2 == 633 || ((pixel_index2 >= 635) && (pixel_index2 <= 637)) || ((pixel_index2 >= 640) && (pixel_index2 <= 643)) || pixel_index2 == 654 || pixel_index2 == 656 || pixel_index2 == 658 || pixel_index2 == 660 || pixel_index2 == 662 || pixel_index2 == 664 || pixel_index2 == 666 || pixel_index2 == 669 || ((pixel_index2 >= 676) && (pixel_index2 <= 677)) || pixel_index2 == 681 || ((pixel_index2 >= 684) && (pixel_index2 <= 685)) || pixel_index2 == 688 || pixel_index2 == 692 || ((pixel_index2 >= 695) && (pixel_index2 <= 696)) || pixel_index2 == 703 || pixel_index2 == 705 || pixel_index2 == 707 || ((pixel_index2 >= 709) && (pixel_index2 <= 710)) || ((pixel_index2 >= 716) && (pixel_index2 <= 717)) || pixel_index2 == 720 || pixel_index2 == 724 || ((pixel_index2 >= 728) && (pixel_index2 <= 729)) || pixel_index2 == 732 || ((pixel_index2 >= 737) && (pixel_index2 <= 739)) || ((pixel_index2 >= 749) && (pixel_index2 <= 750)) || ((pixel_index2 >= 753) && (pixel_index2 <= 754)) || pixel_index2 == 757 || pixel_index2 == 761 || ((pixel_index2 >= 764) && (pixel_index2 <= 765)) || pixel_index2 == 772 || pixel_index2 == 781 || pixel_index2 == 799 || pixel_index2 == 801 || pixel_index2 == 806 || pixel_index2 == 813 || pixel_index2 == 832 || pixel_index2 == 835 || pixel_index2 == 846 || pixel_index2 == 861 || pixel_index2 == 868 || pixel_index2 == 877 || pixel_index2 == 895 || pixel_index2 == 897 || pixel_index2 == 899 || pixel_index2 == 902 || pixel_index2 == 909 || pixel_index2 == 927 || pixel_index2 == 931 || pixel_index2 == 942 || pixel_index2 == 957 || pixel_index2 == 964 || pixel_index2 == 973 || pixel_index2 == 991 || pixel_index2 == 993 || pixel_index2 == 998 || pixel_index2 == 1005 || pixel_index2 == 1023 || pixel_index2 == 1027 || pixel_index2 == 1038 || pixel_index2 == 1052 || ((pixel_index2 >= 1120) && (pixel_index2 <= 1122)) || ((pixel_index2 >= 1634) && (pixel_index2 <= 1635)) || pixel_index2 == 1638 || pixel_index2 == 1640 || pixel_index2 == 1642 || pixel_index2 == 1648 || pixel_index2 == 1651 || pixel_index2 == 1656 || pixel_index2 == 1659 || ((pixel_index2 >= 1665) && (pixel_index2 <= 1666)) || pixel_index2 == 1668 || pixel_index2 == 1672 || pixel_index2 == 1674 || pixel_index2 == 1676 || pixel_index2 == 1678 || ((pixel_index2 >= 1681) && (pixel_index2 <= 1682)) || ((pixel_index2 >= 1686) && (pixel_index2 <= 1687)) || pixel_index2 == 1690 || pixel_index2 == 1692 || ((pixel_index2 >= 1694) && (pixel_index2 <= 1695)) || pixel_index2 == 1700 || pixel_index2 == 1703 || pixel_index2 == 1705 || ((pixel_index2 >= 1707) && (pixel_index2 <= 1708)) || pixel_index2 == 1711 || pixel_index2 == 1715 || ((pixel_index2 >= 1717) && (pixel_index2 <= 1718)) || pixel_index2 == 1721 || ((pixel_index2 >= 1723) && (pixel_index2 <= 1724)) || pixel_index2 == 1732 || pixel_index2 == 1734 || pixel_index2 == 1736 || pixel_index2 == 1739 || pixel_index2 == 1743 || pixel_index2 == 1745 || pixel_index2 == 1748 || pixel_index2 == 1753 || pixel_index2 == 1755 || pixel_index2 == 1760 || pixel_index2 == 1765 || pixel_index2 == 1768 || pixel_index2 == 1770 || pixel_index2 == 1772 || pixel_index2 == 1774 || pixel_index2 == 1776 || pixel_index2 == 1782 || pixel_index2 == 1784 || pixel_index2 == 1786 || pixel_index2 == 1788 || pixel_index2 == 1790 || pixel_index2 == 1792 || pixel_index2 == 1797 || pixel_index2 == 1799 || pixel_index2 == 1801 || pixel_index2 == 1805 || pixel_index2 == 1807 || pixel_index2 == 1809 || pixel_index2 == 1811 || pixel_index2 == 1815 || pixel_index2 == 1817 || pixel_index2 == 1821 || ((pixel_index2 >= 1826) && (pixel_index2 <= 1828)) || pixel_index2 == 1830 || pixel_index2 == 1832 || pixel_index2 == 1835 || pixel_index2 == 1839 || pixel_index2 == 1841 || pixel_index2 == 1844 || pixel_index2 == 1849 || pixel_index2 == 1851 || ((pixel_index2 >= 1857) && (pixel_index2 <= 1858)) || pixel_index2 == 1861 || pixel_index2 == 1864 || pixel_index2 == 1866 || pixel_index2 == 1868 || pixel_index2 == 1870 || ((pixel_index2 >= 1873) && (pixel_index2 <= 1874)) || pixel_index2 == 1878 || pixel_index2 == 1880 || pixel_index2 == 1882 || pixel_index2 == 1884 || pixel_index2 == 1886 || pixel_index2 == 1888 || pixel_index2 == 1893 || pixel_index2 == 1895 || pixel_index2 == 1897 || ((pixel_index2 >= 1899) && (pixel_index2 <= 1901)) || pixel_index2 == 1903 || pixel_index2 == 1905 || pixel_index2 == 1907 || ((pixel_index2 >= 1909) && (pixel_index2 <= 1911)) || pixel_index2 == 1913 || ((pixel_index2 >= 1915) && (pixel_index2 <= 1917)) || pixel_index2 == 1923 || ((pixel_index2 >= 1927) && (pixel_index2 <= 1928)) || ((pixel_index2 >= 1930) && (pixel_index2 <= 1931)) || pixel_index2 == 1936 || ((pixel_index2 >= 1939) && (pixel_index2 <= 1940)) || ((pixel_index2 >= 1944) && (pixel_index2 <= 1945)) || pixel_index2 == 1947 || ((pixel_index2 >= 1952) && (pixel_index2 <= 1953)) || ((pixel_index2 >= 1956) && (pixel_index2 <= 1957)) || ((pixel_index2 >= 1959) && (pixel_index2 <= 1960)) || pixel_index2 == 1962 || ((pixel_index2 >= 1965) && (pixel_index2 <= 1966)) || ((pixel_index2 >= 1968) && (pixel_index2 <= 1969)) || ((pixel_index2 >= 1974) && (pixel_index2 <= 1975)) || ((pixel_index2 >= 1979) && (pixel_index2 <= 1980)) || pixel_index2 == 1983 || ((pixel_index2 >= 1988) && (pixel_index2 <= 1989)) || ((pixel_index2 >= 1992) && (pixel_index2 <= 1993)) || pixel_index2 == 1996 || pixel_index2 == 2000 || ((pixel_index2 >= 2002) && (pixel_index2 <= 2003)) || pixel_index2 == 2006 || pixel_index2 == 2009 || pixel_index2 == 2012 || pixel_index2 == 2024 || pixel_index2 == 2027 || pixel_index2 == 2036 || pixel_index2 == 2041 || pixel_index2 == 2053 || pixel_index2 == 2056 || pixel_index2 == 2062 || pixel_index2 == 2070 || pixel_index2 == 2085 || pixel_index2 == 2105 || pixel_index2 == 2120 || pixel_index2 == 2123 || pixel_index2 == 2132 || pixel_index2 == 2137 || pixel_index2 == 2139 || pixel_index2 == 2149 || pixel_index2 == 2152 || pixel_index2 == 2154 || pixel_index2 == 2158 || pixel_index2 == 2166 || pixel_index2 == 2181 || pixel_index2 == 2201 || pixel_index2 == 2216 || pixel_index2 == 2219 || pixel_index2 == 2228 || pixel_index2 == 2233 || pixel_index2 == 2245 || pixel_index2 == 2247 || pixel_index2 == 2254 || pixel_index2 == 2262 || pixel_index2 == 2277 || pixel_index2 == 2297 || ((pixel_index2 >= 2690) && (pixel_index2 <= 2717)) || ((pixel_index2 >= 2735) && (pixel_index2 <= 2736)) || pixel_index2 == 2830 || pixel_index2 == 2882 || ((pixel_index2 >= 2886) && (pixel_index2 <= 2887)) || ((pixel_index2 >= 2889) && (pixel_index2 <= 2890)) || pixel_index2 == 2893 || pixel_index2 == 2895 || ((pixel_index2 >= 2897) && (pixel_index2 <= 2898)) || pixel_index2 == 2901 || pixel_index2 == 2905 || ((pixel_index2 >= 2908) && (pixel_index2 <= 2909)) || ((pixel_index2 >= 2913) && (pixel_index2 <= 2914)) || pixel_index2 == 2917 || pixel_index2 == 2919 || pixel_index2 == 2921 || pixel_index2 == 2927 || pixel_index2 == 2930 || pixel_index2 == 2932 || pixel_index2 == 2934 || ((pixel_index2 >= 2936) && (pixel_index2 <= 2937)) || pixel_index2 == 2940 || pixel_index2 == 2942 || pixel_index2 == 2944 || pixel_index2 == 2947 || ((pixel_index2 >= 2952) && (pixel_index2 <= 2953)) || pixel_index2 == 2955 || pixel_index2 == 2960 || ((pixel_index2 >= 2962) && (pixel_index2 <= 2963)) || pixel_index2 == 2966 || ((pixel_index2 >= 2970) && (pixel_index2 <= 2972)) || pixel_index2 == 2979 || pixel_index2 == 2981 || pixel_index2 == 2987 || pixel_index2 == 2989 || pixel_index2 == 2991 || pixel_index2 == 2993 || pixel_index2 == 2995 || pixel_index2 == 2997 || pixel_index2 == 2999 || pixel_index2 == 3001 || pixel_index2 == 3003 || pixel_index2 == 3011 || pixel_index2 == 3013 || pixel_index2 == 3015 || pixel_index2 == 3018 || pixel_index2 == 3022 || pixel_index2 == 3024 || pixel_index2 == 3026 || pixel_index2 == 3028 || pixel_index2 == 3030 || pixel_index2 == 3032 || pixel_index2 == 3034 || pixel_index2 == 3036 || pixel_index2 == 3038 || pixel_index2 == 3040 || pixel_index2 == 3043 || pixel_index2 == 3047 || pixel_index2 == 3052 || pixel_index2 == 3056 || pixel_index2 == 3058 || pixel_index2 == 3060 || pixel_index2 == 3063 || pixel_index2 == 3065 || ((pixel_index2 >= 3068) && (pixel_index2 <= 3069)) || pixel_index2 == 3075 || ((pixel_index2 >= 3078) && (pixel_index2 <= 3079)) || ((pixel_index2 >= 3081) && (pixel_index2 <= 3083)) || pixel_index2 == 3085 || pixel_index2 == 3087 || pixel_index2 == 3089 || pixel_index2 == 3091 || pixel_index2 == 3093 || pixel_index2 == 3095 || pixel_index2 == 3097 || ((pixel_index2 >= 3100) && (pixel_index2 <= 3101)) || ((pixel_index2 >= 3105) && (pixel_index2 <= 3107)) || pixel_index2 == 3109 || pixel_index2 == 3111 || pixel_index2 == 3114 || pixel_index2 == 3118 || pixel_index2 == 3120 || pixel_index2 == 3122 || pixel_index2 == 3124 || pixel_index2 == 3126 || pixel_index2 == 3128 || pixel_index2 == 3130 || pixel_index2 == 3132 || pixel_index2 == 3134 || pixel_index2 == 3136 || pixel_index2 == 3139 || ((pixel_index2 >= 3144) && (pixel_index2 <= 3145)) || pixel_index2 == 3148 || pixel_index2 == 3150 || pixel_index2 == 3152 || pixel_index2 == 3154 || pixel_index2 == 3156 || pixel_index2 == 3159 || pixel_index2 == 3161 || ((pixel_index2 >= 3170) && (pixel_index2 <= 3171)) || ((pixel_index2 >= 3173) && (pixel_index2 <= 3174)) || pixel_index2 == 3178 || pixel_index2 == 3181 || pixel_index2 == 3183 || pixel_index2 == 3186 || pixel_index2 == 3190 || ((pixel_index2 >= 3192) && (pixel_index2 <= 3193)) || ((pixel_index2 >= 3195) && (pixel_index2 <= 3196)) || pixel_index2 == 3202 || ((pixel_index2 >= 3206) && (pixel_index2 <= 3207)) || ((pixel_index2 >= 3209) && (pixel_index2 <= 3210)) || ((pixel_index2 >= 3214) && (pixel_index2 <= 3215)) || ((pixel_index2 >= 3219) && (pixel_index2 <= 3220)) || ((pixel_index2 >= 3224) && (pixel_index2 <= 3225)) || ((pixel_index2 >= 3229) && (pixel_index2 <= 3230)) || ((pixel_index2 >= 3234) && (pixel_index2 <= 3235)) || ((pixel_index2 >= 3239) && (pixel_index2 <= 3240)) || ((pixel_index2 >= 3243) && (pixel_index2 <= 3244)) || pixel_index2 == 3247 || pixel_index2 == 3251 || ((pixel_index2 >= 3254) && (pixel_index2 <= 3255)) || ((pixel_index2 >= 3258) && (pixel_index2 <= 3259)) || pixel_index2 == 3267 || pixel_index2 == 3277 || pixel_index2 == 3279 || pixel_index2 == 3303 || pixel_index2 == 3306 || pixel_index2 == 3318 || pixel_index2 == 3320 || pixel_index2 == 3328 || pixel_index2 == 3331 || pixel_index2 == 3340 || pixel_index2 == 3351 || ((pixel_index2 >= 3356) && (pixel_index2 <= 3357)) || pixel_index2 == 3363 || pixel_index2 == 3373 || pixel_index2 == 3375 || pixel_index2 == 3399 || pixel_index2 == 3402 || pixel_index2 == 3416 || pixel_index2 == 3427 || pixel_index2 == 3436 || pixel_index2 == 3447 || pixel_index2 == 3449 || ((pixel_index2 >= 3452) && (pixel_index2 <= 3453)) || pixel_index2 == 3459 || pixel_index2 == 3469 || pixel_index2 == 3471 || pixel_index2 == 3495 || pixel_index2 == 3498 || pixel_index2 == 3512 || pixel_index2 == 3522 || pixel_index2 == 3532 || pixel_index2 == 3543 || ((pixel_index2 >= 3546) && (pixel_index2 <= 3548)) || ((pixel_index2 >= 3840) && (pixel_index2 <= 3936)) || ((pixel_index2 >= 4031) && (pixel_index2 <= 4032)) || ((pixel_index2 >= 4103) && (pixel_index2 <= 4104)) || pixel_index2 == 4110 || ((pixel_index2 >= 4114) && (pixel_index2 <= 4116)) || ((pixel_index2 >= 4120) && (pixel_index2 <= 4123)) || ((pixel_index2 >= 4127) && (pixel_index2 <= 4128)) || pixel_index2 == 4198 || pixel_index2 == 4200 || pixel_index2 == 4206 || pixel_index2 == 4209 || pixel_index2 == 4213 || ((pixel_index2 >= 4215) && (pixel_index2 <= 4216)) || ((pixel_index2 >= 4219) && (pixel_index2 <= 4220)) || ((pixel_index2 >= 4223) && (pixel_index2 <= 4224)) || pixel_index2 == 4296 || pixel_index2 == 4302 || pixel_index2 == 4305 || pixel_index2 == 4309 || ((pixel_index2 >= 4311) && (pixel_index2 <= 4312)) || ((pixel_index2 >= 4319) && (pixel_index2 <= 4320)) || pixel_index2 == 4329 || pixel_index2 == 4392 || pixel_index2 == 4395 || pixel_index2 == 4398 || pixel_index2 == 4401 || pixel_index2 == 4405 || ((pixel_index2 >= 4407) && (pixel_index2 <= 4408)) || ((pixel_index2 >= 4415) && (pixel_index2 <= 4416)) || ((pixel_index2 >= 4424) && (pixel_index2 <= 4426)) || pixel_index2 == 4431 || ((pixel_index2 >= 4486) && (pixel_index2 <= 4489)) || ((pixel_index2 >= 4492) && (pixel_index2 <= 4493)) || pixel_index2 == 4495 || ((pixel_index2 >= 4498) && (pixel_index2 <= 4500)) || ((pixel_index2 >= 4504) && (pixel_index2 <= 4506)) || ((pixel_index2 >= 4511) && (pixel_index2 <= 4512)) || ((pixel_index2 >= 4521) && (pixel_index2 <= 4523)) || ((pixel_index2 >= 4526) && (pixel_index2 <= 4527)) || pixel_index2 == 4584 || ((pixel_index2 >= 4602) && (pixel_index2 <= 4603)) || ((pixel_index2 >= 4607) && (pixel_index2 <= 4608)) || ((pixel_index2 >= 4618) && (pixel_index2 <= 4623)) || pixel_index2 == 4680 || ((pixel_index2 >= 4699) && (pixel_index2 <= 4700)) || ((pixel_index2 >= 4703) && (pixel_index2 <= 4704)) || ((pixel_index2 >= 4715) && (pixel_index2 <= 4720)) || pixel_index2 == 4776 || ((pixel_index2 >= 4791) && (pixel_index2 <= 4792)) || ((pixel_index2 >= 4795) && (pixel_index2 <= 4796)) || ((pixel_index2 >= 4799) && (pixel_index2 <= 4800)) || ((pixel_index2 >= 4811) && (pixel_index2 <= 4816)) || pixel_index2 == 4872 || ((pixel_index2 >= 4888) && (pixel_index2 <= 4891)) || ((pixel_index2 >= 4895) && (pixel_index2 <= 4896)) || ((pixel_index2 >= 4906) && (pixel_index2 <= 4912)) || ((pixel_index2 >= 4991) && (pixel_index2 <= 4992)) || ((pixel_index2 >= 5001) && (pixel_index2 <= 5009)) || ((pixel_index2 >= 5087) && (pixel_index2 <= 5088)) || ((pixel_index2 >= 5099) && (pixel_index2 <= 5105)) || pixel_index2 == 5136 || pixel_index2 == 5140 || ((pixel_index2 >= 5143) && (pixel_index2 <= 5145)) || pixel_index2 == 5148 || ((pixel_index2 >= 5151) && (pixel_index2 <= 5152)) || ((pixel_index2 >= 5156) && (pixel_index2 <= 5158)) || ((pixel_index2 >= 5161) && (pixel_index2 <= 5164)) || pixel_index2 == 5167 || ((pixel_index2 >= 5169) && (pixel_index2 <= 5172)) || ((pixel_index2 >= 5176) && (pixel_index2 <= 5179)) || ((pixel_index2 >= 5183) && (pixel_index2 <= 5184)) || ((pixel_index2 >= 5197) && (pixel_index2 <= 5201)) || pixel_index2 == 5232 || pixel_index2 == 5236 || pixel_index2 == 5238 || pixel_index2 == 5242 || pixel_index2 == 5244 || pixel_index2 == 5246 || pixel_index2 == 5248 || pixel_index2 == 5251 || pixel_index2 == 5255 || pixel_index2 == 5261 || pixel_index2 == 5263 || pixel_index2 == 5269 || ((pixel_index2 >= 5271) && (pixel_index2 <= 5272)) || ((pixel_index2 >= 5275) && (pixel_index2 <= 5276)) || ((pixel_index2 >= 5279) && (pixel_index2 <= 5280)) || ((pixel_index2 >= 5295) && (pixel_index2 <= 5298)) || pixel_index2 == 5328 || pixel_index2 == 5332 || pixel_index2 == 5334 || pixel_index2 == 5338 || pixel_index2 == 5340 || pixel_index2 == 5344 || pixel_index2 == 5351 || ((pixel_index2 >= 5353) && (pixel_index2 <= 5357)) || pixel_index2 == 5359 || ((pixel_index2 >= 5361) && (pixel_index2 <= 5365)) || ((pixel_index2 >= 5367) && (pixel_index2 <= 5368)) || ((pixel_index2 >= 5375) && (pixel_index2 <= 5376)) || ((pixel_index2 >= 5392) && (pixel_index2 <= 5394)) || pixel_index2 == 5424 || pixel_index2 == 5428 || pixel_index2 == 5430 || pixel_index2 == 5434 || pixel_index2 == 5436 || pixel_index2 == 5440 || pixel_index2 == 5443 || pixel_index2 == 5447 || pixel_index2 == 5449 || pixel_index2 == 5453 || pixel_index2 == 5455 || pixel_index2 == 5457 || pixel_index2 == 5461 || ((pixel_index2 >= 5463) && (pixel_index2 <= 5464)) || ((pixel_index2 >= 5471) && (pixel_index2 <= 5472)) || pixel_index2 == 5490 || ((pixel_index2 >= 5521) && (pixel_index2 <= 5524)) || ((pixel_index2 >= 5527) && (pixel_index2 <= 5529)) || pixel_index2 == 5532 || ((pixel_index2 >= 5534) && (pixel_index2 <= 5537)) || ((pixel_index2 >= 5540) && (pixel_index2 <= 5542)) || ((pixel_index2 >= 5546) && (pixel_index2 <= 5548)) || pixel_index2 == 5551 || ((pixel_index2 >= 5554) && (pixel_index2 <= 5556)) || ((pixel_index2 >= 5560) && (pixel_index2 <= 5562)) || ((pixel_index2 >= 5567) && (pixel_index2 <= 5568)) || pixel_index2 == 5632 || pixel_index2 == 5647 || ((pixel_index2 >= 5658) && (pixel_index2 <= 5659)) || ((pixel_index2 >= 5663) && (pixel_index2 <= 5664)) || pixel_index2 == 5724 || pixel_index2 == 5728 || pixel_index2 == 5743 || ((pixel_index2 >= 5755) && (pixel_index2 <= 5756)) || ((pixel_index2 >= 5759) && (pixel_index2 <= 5760)) || pixel_index2 == 5824 || pixel_index2 == 5839 || ((pixel_index2 >= 5847) && (pixel_index2 <= 5848)) || ((pixel_index2 >= 5851) && (pixel_index2 <= 5852)) || ((pixel_index2 >= 5855) && (pixel_index2 <= 5856)) || pixel_index2 == 5920 || pixel_index2 == 5935 || ((pixel_index2 >= 5944) && (pixel_index2 <= 5947)) || ((pixel_index2 >= 5951) && (pixel_index2 <= 5952)) || (pixel_index2 >= 6047) && (pixel_index2 <= 6143)) oled_data2 = 16'b1111011110011110;
        else if (((pixel_index2 >= 4137) && (pixel_index2 <= 4141)) || ((pixel_index2 >= 4153) && (pixel_index2 <= 4157)) || ((pixel_index2 >= 4234) && (pixel_index2 <= 4237)) || ((pixel_index2 >= 4249) && (pixel_index2 <= 4253)) || ((pixel_index2 >= 4331) && (pixel_index2 <= 4333)) || ((pixel_index2 >= 4345) && (pixel_index2 <= 4349)) || ((pixel_index2 >= 4428) && (pixel_index2 <= 4429)) || ((pixel_index2 >= 4441) && (pixel_index2 <= 4445)) || ((pixel_index2 >= 4537) && (pixel_index2 <= 4541)) || ((pixel_index2 >= 4633) && (pixel_index2 <= 4637)) || pixel_index2 == 4713 || ((pixel_index2 >= 4729) && (pixel_index2 <= 4733)) || pixel_index2 == 4809 || ((pixel_index2 >= 4825) && (pixel_index2 <= 4829)) || ((pixel_index2 >= 4921) && (pixel_index2 <= 4925)) || ((pixel_index2 >= 5017) && (pixel_index2 <= 5021)) || ((pixel_index2 >= 5113) && (pixel_index2 <= 5117)) || ((pixel_index2 >= 5193) && (pixel_index2 <= 5194)) || ((pixel_index2 >= 5209) && (pixel_index2 <= 5213)) || ((pixel_index2 >= 5289) && (pixel_index2 <= 5292)) || ((pixel_index2 >= 5305) && (pixel_index2 <= 5309)) || ((pixel_index2 >= 5385) && (pixel_index2 <= 5389)) || (pixel_index2 >= 5481) && (pixel_index2 <= 5485)) oled_data2 = 16'b0000010100000000;
        else oled_data2 = 0;
    end
    else if (sorting_algorithm == 4'b0100) begin //insertion sort
        if (((pixel_index2 >= 0) && (pixel_index2 <= 96)) || ((pixel_index2 >= 191) && (pixel_index2 <= 192)) || ((pixel_index2 >= 287) && (pixel_index2 <= 288)) || ((pixel_index2 >= 383) && (pixel_index2 <= 384)) || ((pixel_index2 >= 479) && (pixel_index2 <= 480)) || ((pixel_index2 >= 575) && (pixel_index2 <= 576)) || ((pixel_index2 >= 671) && (pixel_index2 <= 672)) || ((pixel_index2 >= 767) && (pixel_index2 <= 768)) || ((pixel_index2 >= 863) && (pixel_index2 <= 864)) || ((pixel_index2 >= 959) && (pixel_index2 <= 960)) || ((pixel_index2 >= 1055) && (pixel_index2 <= 1056)) || ((pixel_index2 >= 1151) && (pixel_index2 <= 1152)) || ((pixel_index2 >= 1247) && (pixel_index2 <= 1248)) || ((pixel_index2 >= 1343) && (pixel_index2 <= 1344)) || ((pixel_index2 >= 1439) && (pixel_index2 <= 1440)) || ((pixel_index2 >= 1535) && (pixel_index2 <= 1536)) || ((pixel_index2 >= 1631) && (pixel_index2 <= 1632)) || ((pixel_index2 >= 1727) && (pixel_index2 <= 1728)) || ((pixel_index2 >= 1823) && (pixel_index2 <= 1824)) || ((pixel_index2 >= 1919) && (pixel_index2 <= 1920)) || ((pixel_index2 >= 2015) && (pixel_index2 <= 2016)) || ((pixel_index2 >= 2111) && (pixel_index2 <= 2112)) || ((pixel_index2 >= 2207) && (pixel_index2 <= 2208)) || ((pixel_index2 >= 2303) && (pixel_index2 <= 2304)) || ((pixel_index2 >= 2399) && (pixel_index2 <= 2400)) || ((pixel_index2 >= 2495) && (pixel_index2 <= 2496)) || ((pixel_index2 >= 2591) && (pixel_index2 <= 2592)) || ((pixel_index2 >= 2687) && (pixel_index2 <= 2688)) || ((pixel_index2 >= 2783) && (pixel_index2 <= 2784)) || ((pixel_index2 >= 2879) && (pixel_index2 <= 2880)) || ((pixel_index2 >= 2975) && (pixel_index2 <= 2976)) || ((pixel_index2 >= 3071) && (pixel_index2 <= 3072)) || ((pixel_index2 >= 3167) && (pixel_index2 <= 3168)) || ((pixel_index2 >= 3263) && (pixel_index2 <= 3264)) || ((pixel_index2 >= 3359) && (pixel_index2 <= 3360)) || ((pixel_index2 >= 3455) && (pixel_index2 <= 3456)) || ((pixel_index2 >= 3551) && (pixel_index2 <= 3552)) || ((pixel_index2 >= 3647) && (pixel_index2 <= 3743)) || pixel_index2 == 4149 || pixel_index2 == 4917 || pixel_index2 == 5013 || pixel_index2 == 5105 || pixel_index2 == 5109 || pixel_index2 == 5201 || pixel_index2 == 5205 || pixel_index2 == 5297 || pixel_index2 == 5301 || ((pixel_index2 >= 5393) && (pixel_index2 <= 5394)) || ((pixel_index2 >= 5396) && (pixel_index2 <= 5397)) || ((pixel_index2 >= 5489) && (pixel_index2 <= 5493)) || ((pixel_index2 >= 5585) && (pixel_index2 <= 5589)) || ((pixel_index2 >= 5681) && (pixel_index2 <= 5685)) || (pixel_index2 >= 5777) && (pixel_index2 <= 5781)) oled_data2 = 16'b1111010100000000;
        else if (pixel_index2 == 275 || pixel_index2 == 371 || pixel_index2 == 412 || ((pixel_index2 >= 414) && (pixel_index2 <= 415)) || ((pixel_index2 >= 418) && (pixel_index2 <= 419)) || pixel_index2 == 422 || pixel_index2 == 427 || pixel_index2 == 430 || ((pixel_index2 >= 434) && (pixel_index2 <= 435)) || pixel_index2 == 441 || pixel_index2 == 443 || pixel_index2 == 445 || pixel_index2 == 447 || pixel_index2 == 454 || ((pixel_index2 >= 457) && (pixel_index2 <= 458)) || ((pixel_index2 >= 461) && (pixel_index2 <= 462)) || ((pixel_index2 >= 466) && (pixel_index2 <= 467)) || ((pixel_index2 >= 469) && (pixel_index2 <= 470)) || pixel_index2 == 473 || pixel_index2 == 477 || pixel_index2 == 510 || pixel_index2 == 512 || pixel_index2 == 516 || pixel_index2 == 519 || pixel_index2 == 523 || pixel_index2 == 525 || pixel_index2 == 527 || pixel_index2 == 529 || pixel_index2 == 537 || pixel_index2 == 539 || pixel_index2 == 541 || pixel_index2 == 544 || pixel_index2 == 551 || pixel_index2 == 553 || pixel_index2 == 555 || pixel_index2 == 559 || pixel_index2 == 561 || pixel_index2 == 563 || pixel_index2 == 567 || pixel_index2 == 569 || pixel_index2 == 573 || pixel_index2 == 606 || pixel_index2 == 608 || ((pixel_index2 >= 610) && (pixel_index2 <= 612)) || pixel_index2 == 615 || pixel_index2 == 617 || pixel_index2 == 619 || pixel_index2 == 621 || pixel_index2 == 623 || ((pixel_index2 >= 626) && (pixel_index2 <= 627)) || pixel_index2 == 633 || pixel_index2 == 635 || pixel_index2 == 637 || pixel_index2 == 640 || pixel_index2 == 647 || pixel_index2 == 649 || pixel_index2 == 651 || ((pixel_index2 >= 653) && (pixel_index2 <= 655)) || pixel_index2 == 657 || pixel_index2 == 659 || ((pixel_index2 >= 661) && (pixel_index2 <= 663)) || ((pixel_index2 >= 666) && (pixel_index2 <= 669)) || ((pixel_index2 >= 702) && (pixel_index2 <= 703)) || pixel_index2 == 707 || ((pixel_index2 >= 710) && (pixel_index2 <= 711)) || pixel_index2 == 714 || pixel_index2 == 718 || ((pixel_index2 >= 721) && (pixel_index2 <= 722)) || pixel_index2 == 729 || pixel_index2 == 731 || pixel_index2 == 733 || ((pixel_index2 >= 735) && (pixel_index2 <= 736)) || ((pixel_index2 >= 742) && (pixel_index2 <= 743)) || pixel_index2 == 746 || pixel_index2 == 750 || ((pixel_index2 >= 754) && (pixel_index2 <= 755)) || pixel_index2 == 758 || ((pixel_index2 >= 763) && (pixel_index2 <= 765)) || pixel_index2 == 798 || pixel_index2 == 807 || pixel_index2 == 825 || pixel_index2 == 827 || pixel_index2 == 832 || pixel_index2 == 839 || pixel_index2 == 858 || pixel_index2 == 861 || pixel_index2 == 894 || pixel_index2 == 903 || pixel_index2 == 921 || pixel_index2 == 923 || pixel_index2 == 925 || pixel_index2 == 928 || pixel_index2 == 935 || pixel_index2 == 953 || pixel_index2 == 957 || pixel_index2 == 990 || pixel_index2 == 999 || pixel_index2 == 1017 || pixel_index2 == 1019 || pixel_index2 == 1024 || pixel_index2 == 1031 || pixel_index2 == 1049 || pixel_index2 == 1053 || ((pixel_index2 >= 1146) && (pixel_index2 <= 1148)) || pixel_index2 == 1370 || pixel_index2 == 1398 || pixel_index2 == 1465 || pixel_index2 == 1467 || ((pixel_index2 >= 1493) && (pixel_index2 <= 1495)) || pixel_index2 == 1561 || pixel_index2 == 1590 || pixel_index2 == 1654 || ((pixel_index2 >= 1657) && (pixel_index2 <= 1658)) || pixel_index2 == 1661 || pixel_index2 == 1663 || ((pixel_index2 >= 1665) && (pixel_index2 <= 1666)) || pixel_index2 == 1669 || pixel_index2 == 1671 || pixel_index2 == 1674 || pixel_index2 == 1676 || ((pixel_index2 >= 1678) && (pixel_index2 <= 1679)) || ((pixel_index2 >= 1682) && (pixel_index2 <= 1683)) || ((pixel_index2 >= 1686) && (pixel_index2 <= 1687)) || ((pixel_index2 >= 1690) && (pixel_index2 <= 1691)) || ((pixel_index2 >= 1695) && (pixel_index2 <= 1696)) || pixel_index2 == 1700 || pixel_index2 == 1703 || pixel_index2 == 1705 || ((pixel_index2 >= 1707) && (pixel_index2 <= 1708)) || pixel_index2 == 1711 || pixel_index2 == 1715 || ((pixel_index2 >= 1717) && (pixel_index2 <= 1718)) || pixel_index2 == 1721 || ((pixel_index2 >= 1723) && (pixel_index2 <= 1724)) || pixel_index2 == 1753 || pixel_index2 == 1755 || pixel_index2 == 1757 || pixel_index2 == 1759 || pixel_index2 == 1761 || pixel_index2 == 1763 || pixel_index2 == 1765 || pixel_index2 == 1768 || pixel_index2 == 1770 || pixel_index2 == 1772 || pixel_index2 == 1776 || pixel_index2 == 1778 || pixel_index2 == 1780 || pixel_index2 == 1782 || pixel_index2 == 1784 || pixel_index2 == 1788 || pixel_index2 == 1790 || pixel_index2 == 1797 || pixel_index2 == 1799 || pixel_index2 == 1801 || pixel_index2 == 1805 || pixel_index2 == 1807 || pixel_index2 == 1809 || pixel_index2 == 1811 || pixel_index2 == 1815 || pixel_index2 == 1817 || pixel_index2 == 1821 || pixel_index2 == 1849 || pixel_index2 == 1851 || pixel_index2 == 1853 || pixel_index2 == 1855 || pixel_index2 == 1857 || pixel_index2 == 1859 || pixel_index2 == 1861 || pixel_index2 == 1864 || pixel_index2 == 1866 || pixel_index2 == 1868 || ((pixel_index2 >= 1870) && (pixel_index2 <= 1872)) || pixel_index2 == 1874 || pixel_index2 == 1876 || pixel_index2 == 1878 || pixel_index2 == 1880 || ((pixel_index2 >= 1882) && (pixel_index2 <= 1884)) || ((pixel_index2 >= 1887) && (pixel_index2 <= 1888)) || pixel_index2 == 1893 || pixel_index2 == 1895 || pixel_index2 == 1897 || ((pixel_index2 >= 1899) && (pixel_index2 <= 1901)) || pixel_index2 == 1903 || pixel_index2 == 1905 || pixel_index2 == 1907 || ((pixel_index2 >= 1909) && (pixel_index2 <= 1911)) || pixel_index2 == 1913 || ((pixel_index2 >= 1915) && (pixel_index2 <= 1917)) || pixel_index2 == 1945 || pixel_index2 == 1947 || pixel_index2 == 1949 || pixel_index2 == 1951 || pixel_index2 == 1954 || pixel_index2 == 1957 || ((pixel_index2 >= 1959) && (pixel_index2 <= 1960)) || ((pixel_index2 >= 1963) && (pixel_index2 <= 1964)) || pixel_index2 == 1967 || pixel_index2 == 1970 || pixel_index2 == 1972 || ((pixel_index2 >= 1974) && (pixel_index2 <= 1975)) || pixel_index2 == 1979 || ((pixel_index2 >= 1982) && (pixel_index2 <= 1983)) || ((pixel_index2 >= 1988) && (pixel_index2 <= 1989)) || ((pixel_index2 >= 1992) && (pixel_index2 <= 1993)) || pixel_index2 == 1996 || pixel_index2 == 2000 || ((pixel_index2 >= 2002) && (pixel_index2 <= 2003)) || pixel_index2 == 2006 || pixel_index2 == 2009 || pixel_index2 == 2012 || pixel_index2 == 2045 || pixel_index2 == 2047 || pixel_index2 == 2056 || pixel_index2 == 2085 || pixel_index2 == 2105 || pixel_index2 == 2141 || pixel_index2 == 2143 || pixel_index2 == 2149 || pixel_index2 == 2152 || pixel_index2 == 2181 || pixel_index2 == 2201 || pixel_index2 == 2237 || pixel_index2 == 2239 || pixel_index2 == 2248 || pixel_index2 == 2277 || pixel_index2 == 2297 || ((pixel_index2 >= 2707) && (pixel_index2 <= 2730)) || pixel_index2 == 2766 || pixel_index2 == 2862 || pixel_index2 == 2882 || pixel_index2 == 2884 || pixel_index2 == 2886 || ((pixel_index2 >= 2889) && (pixel_index2 <= 2890)) || ((pixel_index2 >= 2893) && (pixel_index2 <= 2894)) || ((pixel_index2 >= 2900) && (pixel_index2 <= 2901)) || pixel_index2 == 2903 || pixel_index2 == 2908 || ((pixel_index2 >= 2910) && (pixel_index2 <= 2911)) || ((pixel_index2 >= 2915) && (pixel_index2 <= 2916)) || pixel_index2 == 2918 || pixel_index2 == 2920 || pixel_index2 == 2922 || ((pixel_index2 >= 2926) && (pixel_index2 <= 2927)) || pixel_index2 == 2930 || pixel_index2 == 2932 || ((pixel_index2 >= 2934) && (pixel_index2 <= 2935)) || ((pixel_index2 >= 2941) && (pixel_index2 <= 2942)) || ((pixel_index2 >= 2944) && (pixel_index2 <= 2945)) || pixel_index2 == 2950 || ((pixel_index2 >= 2952) && (pixel_index2 <= 2953)) || ((pixel_index2 >= 2957) && (pixel_index2 <= 2958)) || pixel_index2 == 2960 || pixel_index2 == 2964 || pixel_index2 == 2967 || ((pixel_index2 >= 2970) && (pixel_index2 <= 2972)) || pixel_index2 == 2978 || pixel_index2 == 2980 || pixel_index2 == 2983 || pixel_index2 == 2985 || pixel_index2 == 2987 || pixel_index2 == 2991 || pixel_index2 == 2995 || pixel_index2 == 3000 || pixel_index2 == 3004 || pixel_index2 == 3008 || pixel_index2 == 3010 || pixel_index2 == 3014 || pixel_index2 == 3016 || pixel_index2 == 3018 || pixel_index2 == 3022 || pixel_index2 == 3024 || pixel_index2 == 3026 || pixel_index2 == 3028 || pixel_index2 == 3030 || pixel_index2 == 3032 || pixel_index2 == 3036 || pixel_index2 == 3042 || pixel_index2 == 3046 || pixel_index2 == 3048 || pixel_index2 == 3050 || pixel_index2 == 3052 || pixel_index2 == 3054 || pixel_index2 == 3056 || pixel_index2 == 3058 || pixel_index2 == 3060 || pixel_index2 == 3062 || pixel_index2 == 3064 || pixel_index2 == 3066 || pixel_index2 == 3069 || pixel_index2 == 3074 || pixel_index2 == 3076 || pixel_index2 == 3079 || pixel_index2 == 3081 || pixel_index2 == 3083 || ((pixel_index2 >= 3085) && (pixel_index2 <= 3087)) || ((pixel_index2 >= 3092) && (pixel_index2 <= 3093)) || pixel_index2 == 3096 || pixel_index2 == 3098 || pixel_index2 == 3100 || ((pixel_index2 >= 3102) && (pixel_index2 <= 3104)) || ((pixel_index2 >= 3107) && (pixel_index2 <= 3108)) || pixel_index2 == 3110 || pixel_index2 == 3112 || pixel_index2 == 3114 || pixel_index2 == 3118 || pixel_index2 == 3120 || pixel_index2 == 3122 || pixel_index2 == 3124 || pixel_index2 == 3126 || pixel_index2 == 3128 || ((pixel_index2 >= 3133) && (pixel_index2 <= 3134)) || ((pixel_index2 >= 3136) && (pixel_index2 <= 3138)) || pixel_index2 == 3140 || pixel_index2 == 3142 || pixel_index2 == 3144 || pixel_index2 == 3146 || pixel_index2 == 3148 || pixel_index2 == 3150 || pixel_index2 == 3152 || pixel_index2 == 3154 || pixel_index2 == 3156 || pixel_index2 == 3158 || pixel_index2 == 3160 || pixel_index2 == 3165 || ((pixel_index2 >= 3171) && (pixel_index2 <= 3172)) || pixel_index2 == 3174 || pixel_index2 == 3178 || pixel_index2 == 3182 || ((pixel_index2 >= 3187) && (pixel_index2 <= 3188)) || ((pixel_index2 >= 3191) && (pixel_index2 <= 3192)) || pixel_index2 == 3195 || pixel_index2 == 3199 || ((pixel_index2 >= 3202) && (pixel_index2 <= 3203)) || ((pixel_index2 >= 3207) && (pixel_index2 <= 3208)) || pixel_index2 == 3210 || ((pixel_index2 >= 3214) && (pixel_index2 <= 3215)) || ((pixel_index2 >= 3219) && (pixel_index2 <= 3220)) || pixel_index2 == 3223 || ((pixel_index2 >= 3228) && (pixel_index2 <= 3229)) || pixel_index2 == 3233 || pixel_index2 == 3237 || pixel_index2 == 3241 || ((pixel_index2 >= 3245) && (pixel_index2 <= 3246)) || pixel_index2 == 3249 || ((pixel_index2 >= 3251) && (pixel_index2 <= 3252)) || pixel_index2 == 3255 || pixel_index2 == 3261 || pixel_index2 == 3268 || pixel_index2 == 3288 || pixel_index2 == 3310 || pixel_index2 == 3357 || pixel_index2 == 3364 || pixel_index2 == 3384 || pixel_index2 == 3402 || pixel_index2 == 3406 || pixel_index2 == 3450 || pixel_index2 == 3453 || pixel_index2 == 3460 || pixel_index2 == 3480 || pixel_index2 == 3502 || ((pixel_index2 >= 3546) && (pixel_index2 <= 3548)) || ((pixel_index2 >= 3840) && (pixel_index2 <= 3936)) || ((pixel_index2 >= 4031) && (pixel_index2 <= 4032)) || ((pixel_index2 >= 4047) && (pixel_index2 <= 4051)) || ((pixel_index2 >= 4103) && (pixel_index2 <= 4104)) || pixel_index2 == 4110 || ((pixel_index2 >= 4114) && (pixel_index2 <= 4116)) || ((pixel_index2 >= 4120) && (pixel_index2 <= 4123)) || ((pixel_index2 >= 4127) && (pixel_index2 <= 4128)) || ((pixel_index2 >= 4143) && (pixel_index2 <= 4147)) || pixel_index2 == 4198 || pixel_index2 == 4200 || pixel_index2 == 4206 || pixel_index2 == 4209 || pixel_index2 == 4213 || ((pixel_index2 >= 4215) && (pixel_index2 <= 4216)) || ((pixel_index2 >= 4219) && (pixel_index2 <= 4220)) || ((pixel_index2 >= 4223) && (pixel_index2 <= 4224)) || ((pixel_index2 >= 4238) && (pixel_index2 <= 4244)) || pixel_index2 == 4296 || pixel_index2 == 4302 || pixel_index2 == 4305 || pixel_index2 == 4309 || ((pixel_index2 >= 4311) && (pixel_index2 <= 4312)) || ((pixel_index2 >= 4319) && (pixel_index2 <= 4320)) || ((pixel_index2 >= 4334) && (pixel_index2 <= 4340)) || pixel_index2 == 4392 || pixel_index2 == 4395 || pixel_index2 == 4398 || pixel_index2 == 4401 || pixel_index2 == 4405 || ((pixel_index2 >= 4407) && (pixel_index2 <= 4408)) || ((pixel_index2 >= 4415) && (pixel_index2 <= 4416)) || ((pixel_index2 >= 4429) && (pixel_index2 <= 4437)) || ((pixel_index2 >= 4486) && (pixel_index2 <= 4489)) || ((pixel_index2 >= 4492) && (pixel_index2 <= 4493)) || pixel_index2 == 4495 || ((pixel_index2 >= 4498) && (pixel_index2 <= 4500)) || ((pixel_index2 >= 4504) && (pixel_index2 <= 4506)) || ((pixel_index2 >= 4511) && (pixel_index2 <= 4512)) || ((pixel_index2 >= 4525) && (pixel_index2 <= 4533)) || pixel_index2 == 4584 || ((pixel_index2 >= 4602) && (pixel_index2 <= 4603)) || ((pixel_index2 >= 4607) && (pixel_index2 <= 4608)) || ((pixel_index2 >= 4621) && (pixel_index2 <= 4627)) || ((pixel_index2 >= 4629) && (pixel_index2 <= 4630)) || pixel_index2 == 4680 || ((pixel_index2 >= 4699) && (pixel_index2 <= 4700)) || ((pixel_index2 >= 4703) && (pixel_index2 <= 4704)) || pixel_index2 == 4717 || ((pixel_index2 >= 4719) && (pixel_index2 <= 4723)) || pixel_index2 == 4726 || pixel_index2 == 4776 || ((pixel_index2 >= 4791) && (pixel_index2 <= 4792)) || ((pixel_index2 >= 4795) && (pixel_index2 <= 4796)) || ((pixel_index2 >= 4799) && (pixel_index2 <= 4800)) || pixel_index2 == 4813 || pixel_index2 == 4815 || pixel_index2 == 4817 || pixel_index2 == 4819 || pixel_index2 == 4872 || ((pixel_index2 >= 4888) && (pixel_index2 <= 4891)) || ((pixel_index2 >= 4895) && (pixel_index2 <= 4896)) || pixel_index2 == 4911 || pixel_index2 == 4913 || pixel_index2 == 4915 || ((pixel_index2 >= 4991) && (pixel_index2 <= 4992)) || pixel_index2 == 5011 || ((pixel_index2 >= 5087) && (pixel_index2 <= 5088)) || pixel_index2 == 5107 || pixel_index2 == 5132 || pixel_index2 == 5136 || ((pixel_index2 >= 5139) && (pixel_index2 <= 5141)) || pixel_index2 == 5144 || ((pixel_index2 >= 5147) && (pixel_index2 <= 5148)) || pixel_index2 == 5154 || ((pixel_index2 >= 5157) && (pixel_index2 <= 5160)) || ((pixel_index2 >= 5164) && (pixel_index2 <= 5167)) || pixel_index2 == 5169 || pixel_index2 == 5173 || ((pixel_index2 >= 5175) && (pixel_index2 <= 5180)) || ((pixel_index2 >= 5183) && (pixel_index2 <= 5184)) || pixel_index2 == 5203 || pixel_index2 == 5228 || pixel_index2 == 5232 || pixel_index2 == 5234 || pixel_index2 == 5238 || pixel_index2 == 5240 || pixel_index2 == 5242 || pixel_index2 == 5244 || pixel_index2 == 5250 || pixel_index2 == 5257 || pixel_index2 == 5259 || pixel_index2 == 5265 || pixel_index2 == 5269 || ((pixel_index2 >= 5273) && (pixel_index2 <= 5274)) || ((pixel_index2 >= 5279) && (pixel_index2 <= 5280)) || pixel_index2 == 5299 || pixel_index2 == 5324 || pixel_index2 == 5328 || pixel_index2 == 5330 || pixel_index2 == 5334 || pixel_index2 == 5336 || pixel_index2 == 5340 || pixel_index2 == 5346 || ((pixel_index2 >= 5349) && (pixel_index2 <= 5353)) || ((pixel_index2 >= 5356) && (pixel_index2 <= 5358)) || pixel_index2 == 5361 || pixel_index2 == 5365 || ((pixel_index2 >= 5369) && (pixel_index2 <= 5370)) || ((pixel_index2 >= 5375) && (pixel_index2 <= 5376)) || pixel_index2 == 5420 || ((pixel_index2 >= 5423) && (pixel_index2 <= 5424)) || pixel_index2 == 5426 || pixel_index2 == 5430 || pixel_index2 == 5432 || pixel_index2 == 5436 || pixel_index2 == 5439 || pixel_index2 == 5442 || pixel_index2 == 5445 || pixel_index2 == 5449 || pixel_index2 == 5455 || pixel_index2 == 5457 || ((pixel_index2 >= 5460) && (pixel_index2 <= 5461)) || ((pixel_index2 >= 5465) && (pixel_index2 <= 5466)) || ((pixel_index2 >= 5471) && (pixel_index2 <= 5472)) || ((pixel_index2 >= 5517) && (pixel_index2 <= 5518)) || pixel_index2 == 5520 || ((pixel_index2 >= 5523) && (pixel_index2 <= 5525)) || pixel_index2 == 5528 || ((pixel_index2 >= 5530) && (pixel_index2 <= 5533)) || ((pixel_index2 >= 5536) && (pixel_index2 <= 5537)) || pixel_index2 == 5539 || ((pixel_index2 >= 5542) && (pixel_index2 <= 5544)) || ((pixel_index2 >= 5547) && (pixel_index2 <= 5550)) || ((pixel_index2 >= 5554) && (pixel_index2 <= 5555)) || pixel_index2 == 5557 || ((pixel_index2 >= 5561) && (pixel_index2 <= 5562)) || ((pixel_index2 >= 5567) && (pixel_index2 <= 5568)) || pixel_index2 == 5628 || ((pixel_index2 >= 5657) && (pixel_index2 <= 5658)) || ((pixel_index2 >= 5663) && (pixel_index2 <= 5664)) || pixel_index2 == 5720 || pixel_index2 == 5724 || ((pixel_index2 >= 5753) && (pixel_index2 <= 5754)) || ((pixel_index2 >= 5759) && (pixel_index2 <= 5760)) || pixel_index2 == 5820 || ((pixel_index2 >= 5849) && (pixel_index2 <= 5850)) || ((pixel_index2 >= 5855) && (pixel_index2 <= 5856)) || pixel_index2 == 5916 || ((pixel_index2 >= 5943) && (pixel_index2 <= 5948)) || ((pixel_index2 >= 5951) && (pixel_index2 <= 5952)) || (pixel_index2 >= 6047) && (pixel_index2 <= 6143)) oled_data2 = 16'b1111011110011110;
        else if (((pixel_index2 >= 4137) && (pixel_index2 <= 4141)) || ((pixel_index2 >= 4233) && (pixel_index2 <= 4236)) || ((pixel_index2 >= 4329) && (pixel_index2 <= 4332)) || ((pixel_index2 >= 4425) && (pixel_index2 <= 4427)) || ((pixel_index2 >= 4521) && (pixel_index2 <= 4523)) || ((pixel_index2 >= 4617) && (pixel_index2 <= 4619)) || ((pixel_index2 >= 4713) && (pixel_index2 <= 4715)) || ((pixel_index2 >= 4809) && (pixel_index2 <= 4811)) || ((pixel_index2 >= 4905) && (pixel_index2 <= 4908)) || ((pixel_index2 >= 5001) && (pixel_index2 <= 5005)) || ((pixel_index2 >= 5097) && (pixel_index2 <= 5101)) || ((pixel_index2 >= 5193) && (pixel_index2 <= 5197)) || ((pixel_index2 >= 5289) && (pixel_index2 <= 5293)) || ((pixel_index2 >= 5385) && (pixel_index2 <= 5389)) || (pixel_index2 >= 5481) && (pixel_index2 <= 5485)) oled_data2 = 16'b1010000000000000;
        else if (((pixel_index2 >= 4153) && (pixel_index2 <= 4157)) || ((pixel_index2 >= 4249) && (pixel_index2 <= 4253)) || ((pixel_index2 >= 4345) && (pixel_index2 <= 4349)) || ((pixel_index2 >= 4441) && (pixel_index2 <= 4445)) || ((pixel_index2 >= 4537) && (pixel_index2 <= 4541)) || ((pixel_index2 >= 4633) && (pixel_index2 <= 4637)) || ((pixel_index2 >= 4729) && (pixel_index2 <= 4733)) || ((pixel_index2 >= 4825) && (pixel_index2 <= 4829)) || ((pixel_index2 >= 4921) && (pixel_index2 <= 4925)) || ((pixel_index2 >= 5017) && (pixel_index2 <= 5021)) || ((pixel_index2 >= 5113) && (pixel_index2 <= 5117)) || ((pixel_index2 >= 5209) && (pixel_index2 <= 5213)) || (pixel_index2 >= 5305) && (pixel_index2 <= 5309)) oled_data2 = 16'b0000010100000000;
        else oled_data2 = 0;
    end
    else if (sorting_algorithm == 4'b1000) begin //cocktail sort
         // 2nd OLED
         if (pixel_index2 == 0 || ((pixel_index2 >= 95) && (pixel_index2 <= 96)) || ((pixel_index2 >= 191) && (pixel_index2 <= 192)) || ((pixel_index2 >= 287) && (pixel_index2 <= 288)) || ((pixel_index2 >= 383) && (pixel_index2 <= 384)) || ((pixel_index2 >= 479) && (pixel_index2 <= 480)) || ((pixel_index2 >= 575) && (pixel_index2 <= 576)) || ((pixel_index2 >= 671) && (pixel_index2 <= 672)) || ((pixel_index2 >= 767) && (pixel_index2 <= 768)) || ((pixel_index2 >= 863) && (pixel_index2 <= 864)) || ((pixel_index2 >= 959) && (pixel_index2 <= 960)) || ((pixel_index2 >= 1055) && (pixel_index2 <= 1056)) || ((pixel_index2 >= 1151) && (pixel_index2 <= 1152)) || ((pixel_index2 >= 1247) && (pixel_index2 <= 1248)) || ((pixel_index2 >= 1343) && (pixel_index2 <= 1344)) || ((pixel_index2 >= 1439) && (pixel_index2 <= 1440)) || ((pixel_index2 >= 1535) && (pixel_index2 <= 1536)) || ((pixel_index2 >= 1631) && (pixel_index2 <= 1632)) || ((pixel_index2 >= 1727) && (pixel_index2 <= 1728)) || ((pixel_index2 >= 1823) && (pixel_index2 <= 1824)) || ((pixel_index2 >= 1919) && (pixel_index2 <= 1920)) || ((pixel_index2 >= 2015) && (pixel_index2 <= 2016)) || ((pixel_index2 >= 2111) && (pixel_index2 <= 2112)) || ((pixel_index2 >= 2207) && (pixel_index2 <= 2208)) || ((pixel_index2 >= 2303) && (pixel_index2 <= 2304)) || ((pixel_index2 >= 2399) && (pixel_index2 <= 2400)) || ((pixel_index2 >= 2495) && (pixel_index2 <= 2496)) || ((pixel_index2 >= 2591) && (pixel_index2 <= 2592)) || ((pixel_index2 >= 2687) && (pixel_index2 <= 2688)) || ((pixel_index2 >= 2783) && (pixel_index2 <= 2784)) || ((pixel_index2 >= 2879) && (pixel_index2 <= 2880)) || ((pixel_index2 >= 2975) && (pixel_index2 <= 2976)) || ((pixel_index2 >= 3071) && (pixel_index2 <= 3072)) || ((pixel_index2 >= 3167) && (pixel_index2 <= 3168)) || ((pixel_index2 >= 3263) && (pixel_index2 <= 3264)) || ((pixel_index2 >= 3359) && (pixel_index2 <= 3360)) || ((pixel_index2 >= 3455) && (pixel_index2 <= 3456)) || ((pixel_index2 >= 3551) && (pixel_index2 <= 3552)) || ((pixel_index2 >= 3647) && (pixel_index2 <= 3743)) || pixel_index2 == 4727 || pixel_index2 == 4731 || ((pixel_index2 >= 4821) && (pixel_index2 <= 4823)) || pixel_index2 == 4827 || ((pixel_index2 >= 4916) && (pixel_index2 <= 4919)) || pixel_index2 == 4923 || ((pixel_index2 >= 5011) && (pixel_index2 <= 5015)) || ((pixel_index2 >= 5019) && (pixel_index2 <= 5020)) || ((pixel_index2 >= 5107) && (pixel_index2 <= 5111)) || ((pixel_index2 >= 5115) && (pixel_index2 <= 5116)) || pixel_index2 == 5126 || ((pixel_index2 >= 5203) && (pixel_index2 <= 5207)) || ((pixel_index2 >= 5211) && (pixel_index2 <= 5213)) || ((pixel_index2 >= 5222) && (pixel_index2 <= 5224)) || ((pixel_index2 >= 5299) && (pixel_index2 <= 5303)) || ((pixel_index2 >= 5307) && (pixel_index2 <= 5309)) || ((pixel_index2 >= 5318) && (pixel_index2 <= 5319)) || ((pixel_index2 >= 5403) && (pixel_index2 <= 5405)) || (pixel_index2 >= 5499) && (pixel_index2 <= 5502)) oled_data2 = 16'b1111010100000000;
         else if ((pixel_index2 >= 1) && (pixel_index2 <= 94)) oled_data2 = 16'b0101001010000000;
         else if (pixel_index2 == 440 || ((pixel_index2 >= 442) && (pixel_index2 <= 443)) || ((pixel_index2 >= 446) && (pixel_index2 <= 447)) || pixel_index2 == 450 || pixel_index2 == 455 || pixel_index2 == 458 || ((pixel_index2 >= 462) && (pixel_index2 <= 463)) || pixel_index2 == 469 || pixel_index2 == 471 || pixel_index2 == 473 || pixel_index2 == 475 || pixel_index2 == 538 || pixel_index2 == 540 || pixel_index2 == 544 || pixel_index2 == 547 || pixel_index2 == 551 || pixel_index2 == 553 || pixel_index2 == 555 || pixel_index2 == 557 || pixel_index2 == 565 || pixel_index2 == 567 || pixel_index2 == 569 || pixel_index2 == 572 || pixel_index2 == 634 || pixel_index2 == 636 || ((pixel_index2 >= 638) && (pixel_index2 <= 640)) || pixel_index2 == 643 || pixel_index2 == 645 || pixel_index2 == 647 || pixel_index2 == 649 || pixel_index2 == 651 || ((pixel_index2 >= 654) && (pixel_index2 <= 655)) || pixel_index2 == 661 || pixel_index2 == 663 || pixel_index2 == 665 || pixel_index2 == 668 || ((pixel_index2 >= 730) && (pixel_index2 <= 731)) || pixel_index2 == 735 || ((pixel_index2 >= 738) && (pixel_index2 <= 739)) || pixel_index2 == 742 || pixel_index2 == 746 || ((pixel_index2 >= 749) && (pixel_index2 <= 750)) || pixel_index2 == 757 || pixel_index2 == 759 || pixel_index2 == 761 || ((pixel_index2 >= 763) && (pixel_index2 <= 764)) || pixel_index2 == 826 || pixel_index2 == 835 || pixel_index2 == 853 || pixel_index2 == 855 || pixel_index2 == 860 || pixel_index2 == 922 || pixel_index2 == 931 || pixel_index2 == 949 || pixel_index2 == 951 || pixel_index2 == 953 || pixel_index2 == 956 || pixel_index2 == 1018 || pixel_index2 == 1027 || pixel_index2 == 1045 || pixel_index2 == 1047 || pixel_index2 == 1052 || pixel_index2 == 1387 || pixel_index2 == 1482 || pixel_index2 == 1484 || pixel_index2 == 1519 || pixel_index2 == 1578 || pixel_index2 == 1615 || ((pixel_index2 >= 1635) && (pixel_index2 <= 1636)) || pixel_index2 == 1638 || pixel_index2 == 1641 || pixel_index2 == 1643 || ((pixel_index2 >= 1645) && (pixel_index2 <= 1646)) || pixel_index2 == 1649 || pixel_index2 == 1653 || ((pixel_index2 >= 1655) && (pixel_index2 <= 1656)) || pixel_index2 == 1659 || ((pixel_index2 >= 1661) && (pixel_index2 <= 1662)) || ((pixel_index2 >= 1674) && (pixel_index2 <= 1675)) || ((pixel_index2 >= 1679) && (pixel_index2 <= 1680)) || pixel_index2 == 1684 || ((pixel_index2 >= 1686) && (pixel_index2 <= 1687)) || ((pixel_index2 >= 1690) && (pixel_index2 <= 1691)) || pixel_index2 == 1694 || pixel_index2 == 1696 || ((pixel_index2 >= 1706) && (pixel_index2 <= 1707)) || ((pixel_index2 >= 1710) && (pixel_index2 <= 1711)) || ((pixel_index2 >= 1713) && (pixel_index2 <= 1714)) || pixel_index2 == 1718 || pixel_index2 == 1720 || ((pixel_index2 >= 1724) && (pixel_index2 <= 1725)) || pixel_index2 == 1730 || pixel_index2 == 1735 || pixel_index2 == 1737 || pixel_index2 == 1739 || pixel_index2 == 1743 || pixel_index2 == 1745 || pixel_index2 == 1747 || pixel_index2 == 1749 || pixel_index2 == 1753 || pixel_index2 == 1755 || pixel_index2 == 1759 || pixel_index2 == 1770 || pixel_index2 == 1772 || pixel_index2 == 1774 || pixel_index2 == 1776 || pixel_index2 == 1780 || pixel_index2 == 1782 || pixel_index2 == 1784 || pixel_index2 == 1788 || pixel_index2 == 1790 || pixel_index2 == 1792 || pixel_index2 == 1801 || pixel_index2 == 1805 || pixel_index2 == 1807 || pixel_index2 == 1809 || pixel_index2 == 1811 || pixel_index2 == 1813 || pixel_index2 == 1815 || pixel_index2 == 1817 || pixel_index2 == 1819 || ((pixel_index2 >= 1827) && (pixel_index2 <= 1828)) || pixel_index2 == 1831 || pixel_index2 == 1833 || pixel_index2 == 1835 || ((pixel_index2 >= 1837) && (pixel_index2 <= 1839)) || pixel_index2 == 1841 || pixel_index2 == 1843 || pixel_index2 == 1845 || ((pixel_index2 >= 1847) && (pixel_index2 <= 1849)) || pixel_index2 == 1851 || ((pixel_index2 >= 1853) && (pixel_index2 <= 1855)) || pixel_index2 == 1866 || pixel_index2 == 1868 || pixel_index2 == 1870 || pixel_index2 == 1872 || pixel_index2 == 1874 || pixel_index2 == 1876 || pixel_index2 == 1878 || pixel_index2 == 1880 || ((pixel_index2 >= 1882) && (pixel_index2 <= 1884)) || pixel_index2 == 1886 || pixel_index2 == 1888 || ((pixel_index2 >= 1898) && (pixel_index2 <= 1899)) || pixel_index2 == 1901 || pixel_index2 == 1903 || pixel_index2 == 1905 || pixel_index2 == 1907 || pixel_index2 == 1909 || pixel_index2 == 1911 || pixel_index2 == 1913 || ((pixel_index2 >= 1916) && (pixel_index2 <= 1917)) || ((pixel_index2 >= 1922) && (pixel_index2 <= 1923)) || ((pixel_index2 >= 1926) && (pixel_index2 <= 1927)) || ((pixel_index2 >= 1930) && (pixel_index2 <= 1931)) || pixel_index2 == 1934 || pixel_index2 == 1938 || ((pixel_index2 >= 1940) && (pixel_index2 <= 1941)) || pixel_index2 == 1944 || pixel_index2 == 1947 || pixel_index2 == 1950 || pixel_index2 == 1962 || pixel_index2 == 1964 || ((pixel_index2 >= 1967) && (pixel_index2 <= 1968)) || ((pixel_index2 >= 1971) && (pixel_index2 <= 1972)) || pixel_index2 == 1975 || pixel_index2 == 1979 || ((pixel_index2 >= 1983) && (pixel_index2 <= 1984)) || ((pixel_index2 >= 1993) && (pixel_index2 <= 1994)) || ((pixel_index2 >= 1998) && (pixel_index2 <= 1999)) || pixel_index2 == 2002 || pixel_index2 == 2005 || pixel_index2 == 2009 || ((pixel_index2 >= 2011) && (pixel_index2 <= 2012)) || pixel_index2 == 2023 || pixel_index2 == 2043 || pixel_index2 == 2064 || pixel_index2 == 2119 || pixel_index2 == 2139 || pixel_index2 == 2160 || pixel_index2 == 2215 || pixel_index2 == 2235 || pixel_index2 == 2256 || pixel_index2 == 2692 || pixel_index2 == 2787 || pixel_index2 == 2883 || ((pixel_index2 >= 2887) && (pixel_index2 <= 2888)) || pixel_index2 == 2890 || pixel_index2 == 2892 || pixel_index2 == 2895 || pixel_index2 == 2898 || pixel_index2 == 2900 || ((pixel_index2 >= 2903) && (pixel_index2 <= 2904)) || ((pixel_index2 >= 2907) && (pixel_index2 <= 2908)) || pixel_index2 == 2913 || pixel_index2 == 2915 || ((pixel_index2 >= 2917) && (pixel_index2 <= 2918)) || pixel_index2 == 2928 || pixel_index2 == 2930 || pixel_index2 == 2932 || pixel_index2 == 2936 || ((pixel_index2 >= 2940) && (pixel_index2 <= 2941)) || ((pixel_index2 >= 2951) && (pixel_index2 <= 2952)) || ((pixel_index2 >= 2954) && (pixel_index2 <= 2955)) || ((pixel_index2 >= 2959) && (pixel_index2 <= 2960)) || ((pixel_index2 >= 2963) && (pixel_index2 <= 2964)) || ((pixel_index2 >= 2966) && (pixel_index2 <= 2967)) || pixel_index2 == 2973 || pixel_index2 == 2982 || pixel_index2 == 2986 || pixel_index2 == 2988 || pixel_index2 == 2990 || pixel_index2 == 2992 || pixel_index2 == 2994 || pixel_index2 == 2997 || pixel_index2 == 3001 || pixel_index2 == 3005 || pixel_index2 == 3009 || pixel_index2 == 3011 || pixel_index2 == 3013 || pixel_index2 == 3015 || pixel_index2 == 3024 || pixel_index2 == 3026 || pixel_index2 == 3029 || pixel_index2 == 3031 || pixel_index2 == 3033 || pixel_index2 == 3035 || pixel_index2 == 3037 || pixel_index2 == 3046 || pixel_index2 == 3052 || pixel_index2 == 3054 || pixel_index2 == 3058 || pixel_index2 == 3062 || pixel_index2 == 3064 || pixel_index2 == 3069 || ((pixel_index2 >= 3079) && (pixel_index2 <= 3080)) || pixel_index2 == 3082 || pixel_index2 == 3084 || pixel_index2 == 3086 || pixel_index2 == 3088 || pixel_index2 == 3090 || pixel_index2 == 3093 || pixel_index2 == 3097 || ((pixel_index2 >= 3099) && (pixel_index2 <= 3101)) || pixel_index2 == 3103 || pixel_index2 == 3105 || pixel_index2 == 3107 || pixel_index2 == 3109 || pixel_index2 == 3111 || pixel_index2 == 3120 || pixel_index2 == 3122 || pixel_index2 == 3125 || pixel_index2 == 3127 || pixel_index2 == 3129 || pixel_index2 == 3131 || pixel_index2 == 3133 || ((pixel_index2 >= 3143) && (pixel_index2 <= 3144)) || ((pixel_index2 >= 3146) && (pixel_index2 <= 3148)) || ((pixel_index2 >= 3151) && (pixel_index2 <= 3152)) || ((pixel_index2 >= 3155) && (pixel_index2 <= 3156)) || pixel_index2 == 3158 || pixel_index2 == 3160 || pixel_index2 == 3165 || ((pixel_index2 >= 3174) && (pixel_index2 <= 3175)) || ((pixel_index2 >= 3179) && (pixel_index2 <= 3180)) || pixel_index2 == 3183 || pixel_index2 == 3186 || ((pixel_index2 >= 3188) && (pixel_index2 <= 3189)) || ((pixel_index2 >= 3191) && (pixel_index2 <= 3192)) || pixel_index2 == 3196 || ((pixel_index2 >= 3200) && (pixel_index2 <= 3201)) || pixel_index2 == 3203 || ((pixel_index2 >= 3205) && (pixel_index2 <= 3206)) || ((pixel_index2 >= 3217) && (pixel_index2 <= 3218)) || ((pixel_index2 >= 3220) && (pixel_index2 <= 3221)) || pixel_index2 == 3224 || ((pixel_index2 >= 3228) && (pixel_index2 <= 3229)) || ((pixel_index2 >= 3238) && (pixel_index2 <= 3239)) || pixel_index2 == 3243 || ((pixel_index2 >= 3246) && (pixel_index2 <= 3247)) || ((pixel_index2 >= 3250) && (pixel_index2 <= 3251)) || pixel_index2 == 3255 || ((pixel_index2 >= 3259) && (pixel_index2 <= 3261)) || pixel_index2 == 3285 || pixel_index2 == 3301 || pixel_index2 == 3314 || pixel_index2 == 3317 || pixel_index2 == 3325 || pixel_index2 == 3354 || pixel_index2 == 3357 || pixel_index2 == 3378 || pixel_index2 == 3381 || pixel_index2 == 3395 || pixel_index2 == 3397 || pixel_index2 == 3410 || pixel_index2 == 3413 || pixel_index2 == 3421 || pixel_index2 == 3450 || pixel_index2 == 3453 || pixel_index2 == 3477 || pixel_index2 == 3493 || pixel_index2 == 3506 || pixel_index2 == 3509 || pixel_index2 == 3517 || ((pixel_index2 >= 3547) && (pixel_index2 <= 3549)) || ((pixel_index2 >= 3840) && (pixel_index2 <= 3847)) || pixel_index2 == 3849 || ((pixel_index2 >= 3881) && (pixel_index2 <= 3936)) || ((pixel_index2 >= 4031) && (pixel_index2 <= 4032)) || ((pixel_index2 >= 4103) && (pixel_index2 <= 4104)) || pixel_index2 == 4110 || ((pixel_index2 >= 4114) && (pixel_index2 <= 4116)) || ((pixel_index2 >= 4120) && (pixel_index2 <= 4123)) || ((pixel_index2 >= 4127) && (pixel_index2 <= 4128)) || pixel_index2 == 4198 || pixel_index2 == 4200 || pixel_index2 == 4206 || pixel_index2 == 4209 || pixel_index2 == 4213 || ((pixel_index2 >= 4215) && (pixel_index2 <= 4216)) || ((pixel_index2 >= 4219) && (pixel_index2 <= 4220)) || ((pixel_index2 >= 4223) && (pixel_index2 <= 4224)) || pixel_index2 == 4296 || pixel_index2 == 4302 || pixel_index2 == 4305 || pixel_index2 == 4309 || ((pixel_index2 >= 4311) && (pixel_index2 <= 4312)) || ((pixel_index2 >= 4319) && (pixel_index2 <= 4320)) || pixel_index2 == 4392 || pixel_index2 == 4395 || pixel_index2 == 4398 || pixel_index2 == 4401 || pixel_index2 == 4405 || ((pixel_index2 >= 4407) && (pixel_index2 <= 4408)) || ((pixel_index2 >= 4415) && (pixel_index2 <= 4416)) || ((pixel_index2 >= 4486) && (pixel_index2 <= 4489)) || ((pixel_index2 >= 4492) && (pixel_index2 <= 4493)) || pixel_index2 == 4495 || ((pixel_index2 >= 4498) && (pixel_index2 <= 4500)) || ((pixel_index2 >= 4504) && (pixel_index2 <= 4506)) || ((pixel_index2 >= 4511) && (pixel_index2 <= 4512)) || pixel_index2 == 4584 || ((pixel_index2 >= 4602) && (pixel_index2 <= 4603)) || ((pixel_index2 >= 4607) && (pixel_index2 <= 4608)) || pixel_index2 == 4680 || ((pixel_index2 >= 4699) && (pixel_index2 <= 4700)) || ((pixel_index2 >= 4703) && (pixel_index2 <= 4704)) || pixel_index2 == 4776 || ((pixel_index2 >= 4791) && (pixel_index2 <= 4792)) || ((pixel_index2 >= 4795) && (pixel_index2 <= 4796)) || ((pixel_index2 >= 4799) && (pixel_index2 <= 4800)) || pixel_index2 == 4872 || ((pixel_index2 >= 4888) && (pixel_index2 <= 4891)) || ((pixel_index2 >= 4895) && (pixel_index2 <= 4896)) || ((pixel_index2 >= 4991) && (pixel_index2 <= 4992)) || ((pixel_index2 >= 5087) && (pixel_index2 <= 5088)) || pixel_index2 == 5144 || pixel_index2 == 5146 || ((pixel_index2 >= 5148) && (pixel_index2 <= 5151)) || ((pixel_index2 >= 5155) && (pixel_index2 <= 5156)) || pixel_index2 == 5159 || pixel_index2 == 5162 || ((pixel_index2 >= 5165) && (pixel_index2 <= 5166)) || ((pixel_index2 >= 5170) && (pixel_index2 <= 5172)) || ((pixel_index2 >= 5176) && (pixel_index2 <= 5179)) || ((pixel_index2 >= 5183) && (pixel_index2 <= 5184)) || pixel_index2 == 5240 || pixel_index2 == 5242 || pixel_index2 == 5244 || pixel_index2 == 5248 || pixel_index2 == 5250 || pixel_index2 == 5252 || pixel_index2 == 5256 || pixel_index2 == 5258 || pixel_index2 == 5260 || pixel_index2 == 5263 || pixel_index2 == 5265 || pixel_index2 == 5269 || ((pixel_index2 >= 5271) && (pixel_index2 <= 5272)) || ((pixel_index2 >= 5275) && (pixel_index2 <= 5276)) || ((pixel_index2 >= 5279) && (pixel_index2 <= 5280)) || pixel_index2 == 5336 || pixel_index2 == 5338 || pixel_index2 == 5340 || pixel_index2 == 5344 || pixel_index2 == 5348 || ((pixel_index2 >= 5353) && (pixel_index2 <= 5354)) || pixel_index2 == 5359 || pixel_index2 == 5361 || pixel_index2 == 5365 || pixel_index2 == 5372 || ((pixel_index2 >= 5375) && (pixel_index2 <= 5376)) || pixel_index2 == 5432 || pixel_index2 == 5434 || ((pixel_index2 >= 5436) && (pixel_index2 <= 5439)) || pixel_index2 == 5444 || pixel_index2 == 5448 || pixel_index2 == 5450 || pixel_index2 == 5452 || pixel_index2 == 5455 || pixel_index2 == 5457 || pixel_index2 == 5461 || ((pixel_index2 >= 5468) && (pixel_index2 <= 5469)) || ((pixel_index2 >= 5471) && (pixel_index2 <= 5472)) || pixel_index2 == 5528 || pixel_index2 == 5530 || pixel_index2 == 5532 || ((pixel_index2 >= 5538) && (pixel_index2 <= 5541)) || pixel_index2 == 5543 || pixel_index2 == 5546 || ((pixel_index2 >= 5549) && (pixel_index2 <= 5550)) || ((pixel_index2 >= 5554) && (pixel_index2 <= 5556)) || ((pixel_index2 >= 5564) && (pixel_index2 <= 5565)) || ((pixel_index2 >= 5567) && (pixel_index2 <= 5568)) || pixel_index2 == 5624 || ((pixel_index2 >= 5629) && (pixel_index2 <= 5631)) || pixel_index2 == 5636 || pixel_index2 == 5642 || ((pixel_index2 >= 5660) && (pixel_index2 <= 5661)) || ((pixel_index2 >= 5663) && (pixel_index2 <= 5664)) || pixel_index2 == 5720 || pixel_index2 == 5722 || pixel_index2 == 5732 || pixel_index2 == 5738 || pixel_index2 == 5756 || ((pixel_index2 >= 5759) && (pixel_index2 <= 5760)) || pixel_index2 == 5816 || pixel_index2 == 5828 || pixel_index2 == 5834 || ((pixel_index2 >= 5847) && (pixel_index2 <= 5848)) || ((pixel_index2 >= 5851) && (pixel_index2 <= 5852)) || ((pixel_index2 >= 5855) && (pixel_index2 <= 5856)) || pixel_index2 == 5912 || pixel_index2 == 5924 || pixel_index2 == 5930 || ((pixel_index2 >= 5944) && (pixel_index2 <= 5947)) || ((pixel_index2 >= 5951) && (pixel_index2 <= 5952)) || ((pixel_index2 >= 6047) && (pixel_index2 <= 6079)) || ((pixel_index2 >= 6081) && (pixel_index2 <= 6083)) || (pixel_index2 >= 6086) && (pixel_index2 <= 6143)) oled_data2 = 16'b1111011110011110;
         else if (((pixel_index2 >= 3851) && (pixel_index2 <= 3867)) || ((pixel_index2 >= 3947) && (pixel_index2 <= 3962)) || ((pixel_index2 >= 3977) && (pixel_index2 <= 3979)) || ((pixel_index2 >= 4044) && (pixel_index2 <= 4058)) || ((pixel_index2 >= 4073) && (pixel_index2 <= 4075)) || ((pixel_index2 >= 4140) && (pixel_index2 <= 4151)) || ((pixel_index2 >= 4154) && (pixel_index2 <= 4155)) || ((pixel_index2 >= 4169) && (pixel_index2 <= 4171)) || ((pixel_index2 >= 4239) && (pixel_index2 <= 4246)) || ((pixel_index2 >= 4265) && (pixel_index2 <= 4267)) || ((pixel_index2 >= 4336) && (pixel_index2 <= 4343)) || ((pixel_index2 >= 4361) && (pixel_index2 <= 4363)) || ((pixel_index2 >= 4431) && (pixel_index2 <= 4440)) || ((pixel_index2 >= 4456) && (pixel_index2 <= 4459)) || ((pixel_index2 >= 4527) && (pixel_index2 <= 4537)) || ((pixel_index2 >= 4552) && (pixel_index2 <= 4555)) || ((pixel_index2 >= 4627) && (pixel_index2 <= 4630)) || ((pixel_index2 >= 4648) && (pixel_index2 <= 4651)) || ((pixel_index2 >= 4744) && (pixel_index2 <= 4747)) || ((pixel_index2 >= 4841) && (pixel_index2 <= 4843)) || pixel_index2 == 4936 || ((pixel_index2 >= 4938) && (pixel_index2 <= 4939)) || ((pixel_index2 >= 5031) && (pixel_index2 <= 5032)) || ((pixel_index2 >= 5034) && (pixel_index2 <= 5035)) || ((pixel_index2 >= 5130) && (pixel_index2 <= 5131)) || ((pixel_index2 >= 5226) && (pixel_index2 <= 5227)) || ((pixel_index2 >= 5509) && (pixel_index2 <= 5511)) || pixel_index2 == 5600 || ((pixel_index2 >= 5604) && (pixel_index2 <= 5606)) || ((pixel_index2 >= 5695) && (pixel_index2 <= 5702)) || ((pixel_index2 >= 5791) && (pixel_index2 <= 5796)) || pixel_index2 == 5798 || ((pixel_index2 >= 5887) && (pixel_index2 <= 5889)) || ((pixel_index2 >= 5891) && (pixel_index2 <= 5892)) || pixel_index2 == 5984 || pixel_index2 == 5988) oled_data2 = 16'b1010000000000000;
         else if (pixel_index2 == 3872 || pixel_index2 == 3875 || pixel_index2 == 3964 || ((pixel_index2 >= 3968) && (pixel_index2 <= 3969)) || pixel_index2 == 3971 || pixel_index2 == 3974 || pixel_index2 == 4061 || pixel_index2 == 4065 || ((pixel_index2 >= 4070) && (pixel_index2 <= 4071)) || pixel_index2 == 4158 || pixel_index2 == 4162 || ((pixel_index2 >= 4164) && (pixel_index2 <= 4165)) || pixel_index2 == 4167 || ((pixel_index2 >= 4248) && (pixel_index2 <= 4249)) || ((pixel_index2 >= 4254) && (pixel_index2 <= 4256)) || ((pixel_index2 >= 4259) && (pixel_index2 <= 4260)) || pixel_index2 == 4263 || ((pixel_index2 >= 4345) && (pixel_index2 <= 4347)) || pixel_index2 == 4352 || ((pixel_index2 >= 4358) && (pixel_index2 <= 4359)) || pixel_index2 == 4444 || pixel_index2 == 4446 || pixel_index2 == 4450 || pixel_index2 == 4454 || ((pixel_index2 >= 4549) && (pixel_index2 <= 4550)) || ((pixel_index2 >= 4644) && (pixel_index2 <= 4645)) || pixel_index2 == 4741 || pixel_index2 == 4833 || ((pixel_index2 >= 4836) && (pixel_index2 <= 4837)) || pixel_index2 == 4933 || ((pixel_index2 >= 5027) && (pixel_index2 <= 5029)) || pixel_index2 == 5220) oled_data2 = 16'b1010001010000000;
         else if (((pixel_index2 >= 3939) && (pixel_index2 <= 3942)) || ((pixel_index2 >= 4035) && (pixel_index2 <= 4038)) || ((pixel_index2 >= 4131) && (pixel_index2 <= 4135)) || ((pixel_index2 >= 4227) && (pixel_index2 <= 4230)) || ((pixel_index2 >= 4323) && (pixel_index2 <= 4325)) || ((pixel_index2 >= 4332) && (pixel_index2 <= 4333)) || ((pixel_index2 >= 4419) && (pixel_index2 <= 4422)) || ((pixel_index2 >= 4515) && (pixel_index2 <= 4519)) || ((pixel_index2 >= 4611) && (pixel_index2 <= 4615)) || ((pixel_index2 >= 4707) && (pixel_index2 <= 4711)) || ((pixel_index2 >= 4718) && (pixel_index2 <= 4719)) || ((pixel_index2 >= 4803) && (pixel_index2 <= 4807)) || pixel_index2 == 4811 || ((pixel_index2 >= 4813) && (pixel_index2 <= 4815)) || ((pixel_index2 >= 4899) && (pixel_index2 <= 4903)) || ((pixel_index2 >= 4908) && (pixel_index2 <= 4911)) || ((pixel_index2 >= 4995) && (pixel_index2 <= 4999)) || ((pixel_index2 >= 5091) && (pixel_index2 <= 5095)) || ((pixel_index2 >= 5187) && (pixel_index2 <= 5191)) || ((pixel_index2 >= 5283) && (pixel_index2 <= 5287)) || ((pixel_index2 >= 5379) && (pixel_index2 <= 5383)) || ((pixel_index2 >= 5475) && (pixel_index2 <= 5479)) || ((pixel_index2 >= 5571) && (pixel_index2 <= 5575)) || ((pixel_index2 >= 5667) && (pixel_index2 <= 5671)) || ((pixel_index2 >= 5763) && (pixel_index2 <= 5767)) || (pixel_index2 >= 5859) && (pixel_index2 <= 5863)) oled_data2 = 16'b0000010100000000;
         else if (pixel_index2 == 3944 || ((pixel_index2 >= 4040) && (pixel_index2 <= 4042)) || ((pixel_index2 >= 4137) && (pixel_index2 <= 4138)) || ((pixel_index2 >= 4234) && (pixel_index2 <= 4235)) || pixel_index2 == 4327 || pixel_index2 == 4424 || ((pixel_index2 >= 4521) && (pixel_index2 <= 4525)) || ((pixel_index2 >= 4618) && (pixel_index2 <= 4621)) || pixel_index2 == 4716 || ((pixel_index2 >= 4721) && (pixel_index2 <= 4722)) || ((pixel_index2 >= 4817) && (pixel_index2 <= 4819)) || ((pixel_index2 >= 4913) && (pixel_index2 <= 4914)) || pixel_index2 == 5003 || ((pixel_index2 >= 5008) && (pixel_index2 <= 5009)) || ((pixel_index2 >= 5100) && (pixel_index2 <= 5101)) || ((pixel_index2 >= 5104) && (pixel_index2 <= 5105)) || ((pixel_index2 >= 5197) && (pixel_index2 <= 5200)) || ((pixel_index2 >= 5294) && (pixel_index2 <= 5296)) || pixel_index2 == 5391) oled_data2 = 16'b0000000000001010;
         else if (pixel_index2 == 3967 || pixel_index2 == 4060 || pixel_index2 == 4064 || pixel_index2 == 4067 || pixel_index2 == 4069 || pixel_index2 == 4157 || ((pixel_index2 >= 4160) && (pixel_index2 <= 4161)) || pixel_index2 == 4163 || pixel_index2 == 4166 || pixel_index2 == 4253 || ((pixel_index2 >= 4257) && (pixel_index2 <= 4258)) || ((pixel_index2 >= 4261) && (pixel_index2 <= 4262)) || ((pixel_index2 >= 4349) && (pixel_index2 <= 4351)) || ((pixel_index2 >= 4353) && (pixel_index2 <= 4357)) || ((pixel_index2 >= 4442) && (pixel_index2 <= 4443)) || pixel_index2 == 4445 || ((pixel_index2 >= 4447) && (pixel_index2 <= 4449)) || ((pixel_index2 >= 4451) && (pixel_index2 <= 4453)) || ((pixel_index2 >= 4540) && (pixel_index2 <= 4548)) || ((pixel_index2 >= 4636) && (pixel_index2 <= 4643)) || ((pixel_index2 >= 4733) && (pixel_index2 <= 4740)) || ((pixel_index2 >= 4829) && (pixel_index2 <= 4832)) || ((pixel_index2 >= 4834) && (pixel_index2 <= 4835)) || ((pixel_index2 >= 4925) && (pixel_index2 <= 4932)) || ((pixel_index2 >= 5022) && (pixel_index2 <= 5026)) || ((pixel_index2 >= 5118) && (pixel_index2 <= 5124)) || ((pixel_index2 >= 5215) && (pixel_index2 <= 5219)) || ((pixel_index2 >= 5311) && (pixel_index2 <= 5314)) || pixel_index2 == 5316 || ((pixel_index2 >= 5408) && (pixel_index2 <= 5412)) || (pixel_index2 >= 5505) && (pixel_index2 <= 5507)) oled_data2 = 16'b1111001010000000;
         else oled_data2 = 0;
    end
    else if (sorting_algorithm == 4'b0011) begin //celeb
        case (celebframe)
            1: begin
            if (pixel_index2 == 168 || ((pixel_index2 >= 172) && (pixel_index2 <= 175)) || ((pixel_index2 >= 178) && (pixel_index2 <= 180)) || ((pixel_index2 >= 182) && (pixel_index2 <= 185)) || pixel_index2 == 187 || pixel_index2 == 190 || pixel_index2 == 264 || pixel_index2 == 271 || pixel_index2 == 273 || pixel_index2 == 281 || pixel_index2 == 284 || pixel_index2 == 286 || pixel_index2 == 360 || ((pixel_index2 >= 365) && (pixel_index2 <= 367)) || ((pixel_index2 >= 370) && (pixel_index2 <= 371)) || ((pixel_index2 >= 375) && (pixel_index2 <= 377)) || ((pixel_index2 >= 380) && (pixel_index2 <= 382)) || pixel_index2 == 456 || pixel_index2 == 463 || pixel_index2 == 468 || pixel_index2 == 473 || pixel_index2 == 475 || pixel_index2 == 478 || ((pixel_index2 >= 550) && (pixel_index2 <= 554)) || ((pixel_index2 >= 556) && (pixel_index2 <= 559)) || ((pixel_index2 >= 561) && (pixel_index2 <= 563)) || ((pixel_index2 >= 566) && (pixel_index2 <= 569)) || ((pixel_index2 >= 572) && (pixel_index2 <= 574)) || ((pixel_index2 >= 744) && (pixel_index2 <= 746)) || ((pixel_index2 >= 749) && (pixel_index2 <= 751)) || ((pixel_index2 >= 753) && (pixel_index2 <= 756)) || pixel_index2 == 758 || pixel_index2 == 761 || pixel_index2 == 766 || pixel_index2 == 839 || pixel_index2 == 844 || pixel_index2 == 852 || pixel_index2 == 855 || pixel_index2 == 857 || pixel_index2 == 862 || ((pixel_index2 >= 936) && (pixel_index2 <= 937)) || ((pixel_index2 >= 941) && (pixel_index2 <= 942)) || ((pixel_index2 >= 946) && (pixel_index2 <= 948)) || ((pixel_index2 >= 951) && (pixel_index2 <= 953)) || ((pixel_index2 >= 956) && (pixel_index2 <= 958)) || pixel_index2 == 1034 || pixel_index2 == 1039 || pixel_index2 == 1044 || pixel_index2 == 1046 || pixel_index2 == 1049 || pixel_index2 == 1051 || pixel_index2 == 1054 || ((pixel_index2 >= 1127) && (pixel_index2 <= 1129)) || ((pixel_index2 >= 1132) && (pixel_index2 <= 1134)) || ((pixel_index2 >= 1137) && (pixel_index2 <= 1140)) || ((pixel_index2 >= 1143) && (pixel_index2 <= 1145)) || (pixel_index2 >= 1148) && (pixel_index2 <= 1150)) oled_data2 = 16'b1111010100000000;
            else if (pixel_index2 == 2627 || pixel_index2 == 3202 || pixel_index2 == 3392 || pixel_index2 == 3484 || pixel_index2 == 3585 || ((pixel_index2 >= 3674) && (pixel_index2 <= 3675)) || pixel_index2 == 3680 || pixel_index2 == 3773 || ((pixel_index2 >= 3775) && (pixel_index2 <= 3776)) || ((pixel_index2 >= 3867) && (pixel_index2 <= 3869)) || pixel_index2 == 3871 || ((pixel_index2 >= 3962) && (pixel_index2 <= 3964)) || ((pixel_index2 >= 3966) && (pixel_index2 <= 3967)) || ((pixel_index2 >= 4056) && (pixel_index2 <= 4060)) || pixel_index2 == 4062 || ((pixel_index2 >= 4151) && (pixel_index2 <= 4155)) || ((pixel_index2 >= 4246) && (pixel_index2 <= 4250)) || ((pixel_index2 >= 4339) && (pixel_index2 <= 4345)) || pixel_index2 == 4433 || ((pixel_index2 >= 4435) && (pixel_index2 <= 4441)) || ((pixel_index2 >= 4529) && (pixel_index2 <= 4536)) || ((pixel_index2 >= 4624) && (pixel_index2 <= 4631)) || ((pixel_index2 >= 4721) && (pixel_index2 <= 4727)) || ((pixel_index2 >= 4819) && (pixel_index2 <= 4821)) || (pixel_index2 >= 4915) && (pixel_index2 <= 4916)) oled_data2 = 16'b1111001010000000;
            else if (((pixel_index2 >= 4817) && (pixel_index2 <= 4818)) || ((pixel_index2 >= 4911) && (pixel_index2 <= 4914)) || ((pixel_index2 >= 5007) && (pixel_index2 <= 5011)) || ((pixel_index2 >= 5104) && (pixel_index2 <= 5107)) || (pixel_index2 >= 5200) && (pixel_index2 <= 5201)) oled_data2 = 16'b1111011110011110;
            else if (pixel_index2 == 5626 || pixel_index2 == 5630 || ((pixel_index2 >= 5634) && (pixel_index2 <= 5636)) || ((pixel_index2 >= 5638) && (pixel_index2 <= 5641)) || pixel_index2 == 5645 || pixel_index2 == 5649 || pixel_index2 == 5652 || ((pixel_index2 >= 5655) && (pixel_index2 <= 5656)) || ((pixel_index2 >= 5660) && (pixel_index2 <= 5662)) || pixel_index2 == 5729 || pixel_index2 == 5732 || pixel_index2 == 5737 || pixel_index2 == 5741 || pixel_index2 == 5746 || pixel_index2 == 5748 || pixel_index2 == 5750 || pixel_index2 == 5753 || pixel_index2 == 5755 || pixel_index2 == 5818 || pixel_index2 == 5822 || pixel_index2 == 5825 || pixel_index2 == 5828 || ((pixel_index2 >= 5831) && (pixel_index2 <= 5833)) || pixel_index2 == 5837 || ((pixel_index2 >= 5842) && (pixel_index2 <= 5844)) || pixel_index2 == 5846 || pixel_index2 == 5849 || ((pixel_index2 >= 5852) && (pixel_index2 <= 5853)) || pixel_index2 == 5914 || pixel_index2 == 5918 || pixel_index2 == 5921 || pixel_index2 == 5924 || pixel_index2 == 5929 || pixel_index2 == 5933 || pixel_index2 == 5937 || pixel_index2 == 5940 || pixel_index2 == 5942 || pixel_index2 == 5945 || pixel_index2 == 5950 || pixel_index2 == 6010 || pixel_index2 == 6014 || ((pixel_index2 >= 6018) && (pixel_index2 <= 6020)) || ((pixel_index2 >= 6022) && (pixel_index2 <= 6025)) || ((pixel_index2 >= 6027) && (pixel_index2 <= 6031)) || ((pixel_index2 >= 6034) && (pixel_index2 <= 6036)) || ((pixel_index2 >= 6039) && (pixel_index2 <= 6040)) || (pixel_index2 >= 6043) && (pixel_index2 <= 6045)) oled_data2 = 16'b0000010100000000;
            else oled_data2 = 0;
            end
            2: begin
            if (pixel_index2 == 168 || ((pixel_index2 >= 172) && (pixel_index2 <= 175)) || ((pixel_index2 >= 178) && (pixel_index2 <= 180)) || ((pixel_index2 >= 182) && (pixel_index2 <= 185)) || pixel_index2 == 187 || pixel_index2 == 190 || pixel_index2 == 264 || pixel_index2 == 271 || pixel_index2 == 273 || pixel_index2 == 281 || pixel_index2 == 284 || pixel_index2 == 286 || pixel_index2 == 360 || ((pixel_index2 >= 365) && (pixel_index2 <= 367)) || ((pixel_index2 >= 370) && (pixel_index2 <= 371)) || ((pixel_index2 >= 375) && (pixel_index2 <= 377)) || ((pixel_index2 >= 380) && (pixel_index2 <= 382)) || pixel_index2 == 456 || pixel_index2 == 463 || pixel_index2 == 468 || pixel_index2 == 473 || pixel_index2 == 475 || pixel_index2 == 478 || ((pixel_index2 >= 550) && (pixel_index2 <= 554)) || ((pixel_index2 >= 556) && (pixel_index2 <= 559)) || ((pixel_index2 >= 561) && (pixel_index2 <= 563)) || ((pixel_index2 >= 566) && (pixel_index2 <= 569)) || ((pixel_index2 >= 572) && (pixel_index2 <= 574)) || ((pixel_index2 >= 744) && (pixel_index2 <= 746)) || ((pixel_index2 >= 749) && (pixel_index2 <= 751)) || ((pixel_index2 >= 753) && (pixel_index2 <= 756)) || pixel_index2 == 758 || pixel_index2 == 761 || pixel_index2 == 766 || pixel_index2 == 839 || pixel_index2 == 844 || pixel_index2 == 852 || pixel_index2 == 855 || pixel_index2 == 857 || pixel_index2 == 862 || ((pixel_index2 >= 936) && (pixel_index2 <= 937)) || ((pixel_index2 >= 941) && (pixel_index2 <= 942)) || ((pixel_index2 >= 946) && (pixel_index2 <= 948)) || ((pixel_index2 >= 951) && (pixel_index2 <= 953)) || ((pixel_index2 >= 956) && (pixel_index2 <= 958)) || pixel_index2 == 1034 || pixel_index2 == 1039 || pixel_index2 == 1044 || pixel_index2 == 1046 || pixel_index2 == 1049 || pixel_index2 == 1051 || pixel_index2 == 1054 || ((pixel_index2 >= 1127) && (pixel_index2 <= 1129)) || ((pixel_index2 >= 1132) && (pixel_index2 <= 1134)) || ((pixel_index2 >= 1137) && (pixel_index2 <= 1140)) || ((pixel_index2 >= 1143) && (pixel_index2 <= 1145)) || (pixel_index2 >= 1148) && (pixel_index2 <= 1150)) oled_data2 = 16'b1111000000001010;
            else if (((pixel_index2 >= 3581) && (pixel_index2 <= 3582)) || ((pixel_index2 >= 3663) && (pixel_index2 <= 3664)) || ((pixel_index2 >= 3670) && (pixel_index2 <= 3671)) || ((pixel_index2 >= 3677) && (pixel_index2 <= 3678)) || ((pixel_index2 >= 3759) && (pixel_index2 <= 3760)) || ((pixel_index2 >= 3766) && (pixel_index2 <= 3767)) || ((pixel_index2 >= 3845) && (pixel_index2 <= 3846)) || ((pixel_index2 >= 3874) && (pixel_index2 <= 3875)) || ((pixel_index2 >= 3941) && (pixel_index2 <= 3942)) || ((pixel_index2 >= 3970) && (pixel_index2 <= 3971)) || ((pixel_index2 >= 4224) && (pixel_index2 <= 4225)) || ((pixel_index2 >= 4320) && (pixel_index2 <= 4321)) || pixel_index2 == 4818 || ((pixel_index2 >= 4839) && (pixel_index2 <= 4840)) || ((pixel_index2 >= 4896) && (pixel_index2 <= 4897)) || ((pixel_index2 >= 4913) && (pixel_index2 <= 4914)) || ((pixel_index2 >= 4935) && (pixel_index2 <= 4936)) || ((pixel_index2 >= 4992) && (pixel_index2 <= 4993)) || ((pixel_index2 >= 5008) && (pixel_index2 <= 5012)) || ((pixel_index2 >= 5103) && (pixel_index2 <= 5107)) || pixel_index2 == 5201 || ((pixel_index2 >= 5203) && (pixel_index2 <= 5204)) || ((pixel_index2 >= 5571) && (pixel_index2 <= 5572)) || ((pixel_index2 >= 5667) && (pixel_index2 <= 5668)) || (pixel_index2 >= 6065) && (pixel_index2 <= 6066)) oled_data2 = 16'b1111011110011110;
            else if (pixel_index2 == 3773 || pixel_index2 == 3857 || pixel_index2 == 3862 || ((pixel_index2 >= 3868) && (pixel_index2 <= 3869)) || pixel_index2 == 3947 || pixel_index2 == 3953 || pixel_index2 == 3958 || pixel_index2 == 3964 || pixel_index2 == 4038 || pixel_index2 == 4043 || pixel_index2 == 4049 || ((pixel_index2 >= 4053) && (pixel_index2 <= 4054)) || ((pixel_index2 >= 4059) && (pixel_index2 <= 4060)) || pixel_index2 == 4066 || pixel_index2 == 4132 || ((pixel_index2 >= 4134) && (pixel_index2 <= 4135)) || ((pixel_index2 >= 4139) && (pixel_index2 <= 4140)) || pixel_index2 == 4149 || pixel_index2 == 4155 || pixel_index2 == 4158 || ((pixel_index2 >= 4161) && (pixel_index2 <= 4162)) || pixel_index2 == 4229 || ((pixel_index2 >= 4231) && (pixel_index2 <= 4233)) || pixel_index2 == 4236 || pixel_index2 == 4244 || pixel_index2 == 4250 || ((pixel_index2 >= 4253) && (pixel_index2 <= 4254)) || pixel_index2 == 4257 || pixel_index2 == 4322 || pixel_index2 == 4325 || ((pixel_index2 >= 4329) && (pixel_index2 <= 4335)) || pixel_index2 == 4340 || ((pixel_index2 >= 4344) && (pixel_index2 <= 4345)) || pixel_index2 == 4349 || pixel_index2 == 4353 || pixel_index2 == 4419 || ((pixel_index2 >= 4429) && (pixel_index2 <= 4430)) || ((pixel_index2 >= 4435) && (pixel_index2 <= 4436)) || ((pixel_index2 >= 4438) && (pixel_index2 <= 4441)) || ((pixel_index2 >= 4443) && (pixel_index2 <= 4444)) || ((pixel_index2 >= 4448) && (pixel_index2 <= 4449)) || pixel_index2 == 4516 || pixel_index2 == 4523 || pixel_index2 == 4526 || pixel_index2 == 4535 || pixel_index2 == 4544 || ((pixel_index2 >= 4615) && (pixel_index2 <= 4617)) || ((pixel_index2 >= 4622) && (pixel_index2 <= 4623)) || ((pixel_index2 >= 4628) && (pixel_index2 <= 4629)) || pixel_index2 == 4631 || pixel_index2 == 4708 || ((pixel_index2 >= 4716) && (pixel_index2 <= 4717)) || pixel_index2 == 4720 || ((pixel_index2 >= 4723) && (pixel_index2 <= 4724)) || pixel_index2 == 4726 || ((pixel_index2 >= 4729) && (pixel_index2 <= 4730)) || ((pixel_index2 >= 4732) && (pixel_index2 <= 4733)) || pixel_index2 == 4738 || ((pixel_index2 >= 4804) && (pixel_index2 <= 4805)) || pixel_index2 == 4810 || pixel_index2 == 4822 || pixel_index2 == 4825 || pixel_index2 == 4828 || ((pixel_index2 >= 4833) && (pixel_index2 <= 4834)) || pixel_index2 == 4898 || ((pixel_index2 >= 4901) && (pixel_index2 <= 4902)) || ((pixel_index2 >= 4907) && (pixel_index2 <= 4908)) || ((pixel_index2 >= 4920) && (pixel_index2 <= 4923)) || ((pixel_index2 >= 4928) && (pixel_index2 <= 4929)) || pixel_index2 == 4934 || ((pixel_index2 >= 4994) && (pixel_index2 <= 4996)) || ((pixel_index2 >= 4998) && (pixel_index2 <= 4999)) || pixel_index2 == 5001 || ((pixel_index2 >= 5004) && (pixel_index2 <= 5005)) || ((pixel_index2 >= 5017) && (pixel_index2 <= 5018)) || ((pixel_index2 >= 5022) && (pixel_index2 <= 5023)) || pixel_index2 == 5029 || ((pixel_index2 >= 5111) && (pixel_index2 <= 5113)) || pixel_index2 == 5116 || ((pixel_index2 >= 5123) && (pixel_index2 <= 5124)) || pixel_index2 == 5195 || ((pixel_index2 >= 5217) && (pixel_index2 <= 5218)) || ((pixel_index2 >= 5285) && (pixel_index2 <= 5286)) || ((pixel_index2 >= 5290) && (pixel_index2 <= 5293)) || ((pixel_index2 >= 5312) && (pixel_index2 <= 5313)) || ((pixel_index2 >= 5382) && (pixel_index2 <= 5384)) || ((pixel_index2 >= 5392) && (pixel_index2 <= 5394)) || pixel_index2 == 5485 || pixel_index2 == 5487 || pixel_index2 == 5491 || pixel_index2 == 5503 || ((pixel_index2 >= 5573) && (pixel_index2 <= 5574)) || pixel_index2 == 5581 || pixel_index2 == 5585 || pixel_index2 == 5588 || ((pixel_index2 >= 5590) && (pixel_index2 <= 5591)) || ((pixel_index2 >= 5598) && (pixel_index2 <= 5599)) || pixel_index2 == 5626 || pixel_index2 == 5630 || ((pixel_index2 >= 5634) && (pixel_index2 <= 5636)) || ((pixel_index2 >= 5638) && (pixel_index2 <= 5641)) || pixel_index2 == 5645 || pixel_index2 == 5649 || pixel_index2 == 5652 || ((pixel_index2 >= 5655) && (pixel_index2 <= 5656)) || ((pixel_index2 >= 5660) && (pixel_index2 <= 5662)) || ((pixel_index2 >= 5684) && (pixel_index2 <= 5689)) || ((pixel_index2 >= 5692) && (pixel_index2 <= 5693)) || pixel_index2 == 5729 || pixel_index2 == 5732 || pixel_index2 == 5737 || pixel_index2 == 5741 || pixel_index2 == 5746 || pixel_index2 == 5748 || pixel_index2 == 5750 || pixel_index2 == 5753 || pixel_index2 == 5755 || pixel_index2 == 5777 || ((pixel_index2 >= 5785) && (pixel_index2 <= 5787)) || pixel_index2 == 5818 || pixel_index2 == 5822 || pixel_index2 == 5825 || pixel_index2 == 5828 || ((pixel_index2 >= 5831) && (pixel_index2 <= 5833)) || pixel_index2 == 5837 || ((pixel_index2 >= 5842) && (pixel_index2 <= 5844)) || pixel_index2 == 5846 || pixel_index2 == 5849 || ((pixel_index2 >= 5852) && (pixel_index2 <= 5853)) || pixel_index2 == 5873 || pixel_index2 == 5914 || pixel_index2 == 5918 || pixel_index2 == 5921 || pixel_index2 == 5924 || pixel_index2 == 5929 || pixel_index2 == 5933 || pixel_index2 == 5937 || pixel_index2 == 5940 || pixel_index2 == 5942 || pixel_index2 == 5945 || pixel_index2 == 5950 || pixel_index2 == 5969 || pixel_index2 == 6010 || pixel_index2 == 6014 || ((pixel_index2 >= 6018) && (pixel_index2 <= 6020)) || ((pixel_index2 >= 6022) && (pixel_index2 <= 6025)) || ((pixel_index2 >= 6027) && (pixel_index2 <= 6031)) || ((pixel_index2 >= 6034) && (pixel_index2 <= 6036)) || ((pixel_index2 >= 6039) && (pixel_index2 <= 6040)) || (pixel_index2 >= 6043) && (pixel_index2 <= 6045)) oled_data2 = 16'b1010000000000000;
            else if (pixel_index2 == 4241 || pixel_index2 == 4337 || pixel_index2 == 4433 || pixel_index2 == 4529 || pixel_index2 == 4534 || ((pixel_index2 >= 4625) && (pixel_index2 <= 4626)) || pixel_index2 == 4630 || ((pixel_index2 >= 4713) && (pixel_index2 <= 4715)) || ((pixel_index2 >= 4718) && (pixel_index2 <= 4719)) || ((pixel_index2 >= 4721) && (pixel_index2 <= 4722)) || pixel_index2 == 4725 || pixel_index2 == 4728 || ((pixel_index2 >= 4811) && (pixel_index2 <= 4817)) || ((pixel_index2 >= 4819) && (pixel_index2 <= 4821)) || ((pixel_index2 >= 4823) && (pixel_index2 <= 4824)) || ((pixel_index2 >= 4909) && (pixel_index2 <= 4912)) || ((pixel_index2 >= 4915) && (pixel_index2 <= 4919)) || ((pixel_index2 >= 5002) && (pixel_index2 <= 5003)) || ((pixel_index2 >= 5006) && (pixel_index2 <= 5007)) || ((pixel_index2 >= 5013) && (pixel_index2 <= 5016)) || ((pixel_index2 >= 5098) && (pixel_index2 <= 5102)) || ((pixel_index2 >= 5108) && (pixel_index2 <= 5110)) || ((pixel_index2 >= 5196) && (pixel_index2 <= 5200)) || pixel_index2 == 5202 || pixel_index2 == 5205 || ((pixel_index2 >= 5294) && (pixel_index2 <= 5302)) || ((pixel_index2 >= 5390) && (pixel_index2 <= 5391)) || ((pixel_index2 >= 5395) && (pixel_index2 <= 5400)) || pixel_index2 == 5486 || ((pixel_index2 >= 5492) && (pixel_index2 <= 5497)) || pixel_index2 == 5582 || pixel_index2 == 5589) oled_data2 = 16'b1111010100010100;
            else oled_data2 = 0;
            end
            3: begin
            if (((pixel_index2 >= 66) && (pixel_index2 <= 69)) || ((pixel_index2 >= 161) && (pixel_index2 <= 165)) || ((pixel_index2 >= 257) && (pixel_index2 <= 261)) || ((pixel_index2 >= 353) && (pixel_index2 <= 357)) || ((pixel_index2 >= 450) && (pixel_index2 <= 453)) || ((pixel_index2 >= 545) && (pixel_index2 <= 549)) || ((pixel_index2 >= 641) && (pixel_index2 <= 646)) || ((pixel_index2 >= 738) && (pixel_index2 <= 742)) || ((pixel_index2 >= 834) && (pixel_index2 <= 836)) || pixel_index2 == 838 || (pixel_index2 >= 930) && (pixel_index2 <= 932)) oled_data2 = 16'b1111001010000000;
            else if (pixel_index2 == 168 || ((pixel_index2 >= 172) && (pixel_index2 <= 175)) || ((pixel_index2 >= 178) && (pixel_index2 <= 180)) || ((pixel_index2 >= 182) && (pixel_index2 <= 185)) || pixel_index2 == 187 || pixel_index2 == 190 || pixel_index2 == 264 || pixel_index2 == 271 || pixel_index2 == 273 || pixel_index2 == 281 || pixel_index2 == 284 || pixel_index2 == 286 || pixel_index2 == 360 || ((pixel_index2 >= 365) && (pixel_index2 <= 367)) || ((pixel_index2 >= 370) && (pixel_index2 <= 371)) || ((pixel_index2 >= 375) && (pixel_index2 <= 377)) || ((pixel_index2 >= 380) && (pixel_index2 <= 382)) || pixel_index2 == 456 || pixel_index2 == 463 || pixel_index2 == 468 || pixel_index2 == 473 || pixel_index2 == 475 || pixel_index2 == 478 || ((pixel_index2 >= 550) && (pixel_index2 <= 554)) || ((pixel_index2 >= 556) && (pixel_index2 <= 559)) || ((pixel_index2 >= 561) && (pixel_index2 <= 563)) || ((pixel_index2 >= 566) && (pixel_index2 <= 569)) || ((pixel_index2 >= 572) && (pixel_index2 <= 574)) || ((pixel_index2 >= 744) && (pixel_index2 <= 746)) || ((pixel_index2 >= 749) && (pixel_index2 <= 751)) || ((pixel_index2 >= 753) && (pixel_index2 <= 756)) || pixel_index2 == 758 || pixel_index2 == 761 || pixel_index2 == 766 || pixel_index2 == 839 || pixel_index2 == 844 || pixel_index2 == 852 || pixel_index2 == 855 || pixel_index2 == 857 || pixel_index2 == 862 || ((pixel_index2 >= 936) && (pixel_index2 <= 937)) || ((pixel_index2 >= 941) && (pixel_index2 <= 942)) || ((pixel_index2 >= 946) && (pixel_index2 <= 948)) || ((pixel_index2 >= 951) && (pixel_index2 <= 953)) || ((pixel_index2 >= 956) && (pixel_index2 <= 958)) || pixel_index2 == 1034 || pixel_index2 == 1039 || pixel_index2 == 1044 || pixel_index2 == 1046 || pixel_index2 == 1049 || pixel_index2 == 1051 || pixel_index2 == 1054 || ((pixel_index2 >= 1127) && (pixel_index2 <= 1129)) || ((pixel_index2 >= 1132) && (pixel_index2 <= 1134)) || ((pixel_index2 >= 1137) && (pixel_index2 <= 1140)) || ((pixel_index2 >= 1143) && (pixel_index2 <= 1145)) || (pixel_index2 >= 1148) && (pixel_index2 <= 1150)) oled_data2 = 16'b0000011110011110;
            else if (pixel_index2 == 837 || ((pixel_index2 >= 933) && (pixel_index2 <= 935)) || ((pixel_index2 >= 1028) && (pixel_index2 <= 1031)) || ((pixel_index2 >= 1124) && (pixel_index2 <= 1126)) || ((pixel_index2 >= 1221) && (pixel_index2 <= 1223)) || ((pixel_index2 >= 3581) && (pixel_index2 <= 3582)) || ((pixel_index2 >= 3663) && (pixel_index2 <= 3664)) || ((pixel_index2 >= 3670) && (pixel_index2 <= 3671)) || ((pixel_index2 >= 3677) && (pixel_index2 <= 3678)) || ((pixel_index2 >= 3759) && (pixel_index2 <= 3760)) || ((pixel_index2 >= 3766) && (pixel_index2 <= 3767)) || ((pixel_index2 >= 3845) && (pixel_index2 <= 3846)) || ((pixel_index2 >= 3874) && (pixel_index2 <= 3875)) || ((pixel_index2 >= 3941) && (pixel_index2 <= 3942)) || ((pixel_index2 >= 3970) && (pixel_index2 <= 3971)) || ((pixel_index2 >= 4224) && (pixel_index2 <= 4225)) || ((pixel_index2 >= 4320) && (pixel_index2 <= 4321)) || ((pixel_index2 >= 4839) && (pixel_index2 <= 4840)) || ((pixel_index2 >= 4896) && (pixel_index2 <= 4897)) || ((pixel_index2 >= 4935) && (pixel_index2 <= 4936)) || ((pixel_index2 >= 4992) && (pixel_index2 <= 4993)) || ((pixel_index2 >= 5571) && (pixel_index2 <= 5572)) || ((pixel_index2 >= 5667) && (pixel_index2 <= 5668)) || (pixel_index2 >= 6065) && (pixel_index2 <= 6066)) oled_data2 = 16'b1111011110011110;
            else if (pixel_index2 == 3773 || pixel_index2 == 3857 || pixel_index2 == 3862 || ((pixel_index2 >= 3868) && (pixel_index2 <= 3869)) || pixel_index2 == 3947 || pixel_index2 == 3953 || pixel_index2 == 3958 || pixel_index2 == 3964 || pixel_index2 == 4038 || pixel_index2 == 4043 || pixel_index2 == 4049 || ((pixel_index2 >= 4053) && (pixel_index2 <= 4054)) || ((pixel_index2 >= 4059) && (pixel_index2 <= 4060)) || pixel_index2 == 4066 || pixel_index2 == 4132 || ((pixel_index2 >= 4134) && (pixel_index2 <= 4135)) || ((pixel_index2 >= 4139) && (pixel_index2 <= 4140)) || ((pixel_index2 >= 4145) && (pixel_index2 <= 4146)) || pixel_index2 == 4149 || pixel_index2 == 4155 || pixel_index2 == 4158 || ((pixel_index2 >= 4161) && (pixel_index2 <= 4162)) || pixel_index2 == 4229 || ((pixel_index2 >= 4231) && (pixel_index2 <= 4233)) || pixel_index2 == 4236 || ((pixel_index2 >= 4241) && (pixel_index2 <= 4242)) || pixel_index2 == 4244 || ((pixel_index2 >= 4249) && (pixel_index2 <= 4251)) || ((pixel_index2 >= 4253) && (pixel_index2 <= 4254)) || pixel_index2 == 4257 || pixel_index2 == 4322 || pixel_index2 == 4325 || ((pixel_index2 >= 4329) && (pixel_index2 <= 4333)) || ((pixel_index2 >= 4337) && (pixel_index2 <= 4338)) || ((pixel_index2 >= 4340) && (pixel_index2 <= 4341)) || ((pixel_index2 >= 4345) && (pixel_index2 <= 4347)) || pixel_index2 == 4349 || pixel_index2 == 4353 || pixel_index2 == 4419 || ((pixel_index2 >= 4427) && (pixel_index2 <= 4430)) || ((pixel_index2 >= 4433) && (pixel_index2 <= 4437)) || ((pixel_index2 >= 4442) && (pixel_index2 <= 4444)) || ((pixel_index2 >= 4448) && (pixel_index2 <= 4449)) || pixel_index2 == 4516 || ((pixel_index2 >= 4523) && (pixel_index2 <= 4526)) || ((pixel_index2 >= 4531) && (pixel_index2 <= 4532)) || ((pixel_index2 >= 4538) && (pixel_index2 <= 4539)) || pixel_index2 == 4544 || ((pixel_index2 >= 4615) && (pixel_index2 <= 4617)) || ((pixel_index2 >= 4634) && (pixel_index2 <= 4635)) || pixel_index2 == 4708 || pixel_index2 == 4713 || ((pixel_index2 >= 4732) && (pixel_index2 <= 4733)) || pixel_index2 == 4738 || ((pixel_index2 >= 4804) && (pixel_index2 <= 4805)) || ((pixel_index2 >= 4833) && (pixel_index2 <= 4834)) || pixel_index2 == 4898 || ((pixel_index2 >= 4901) && (pixel_index2 <= 4902)) || ((pixel_index2 >= 4928) && (pixel_index2 <= 4929)) || pixel_index2 == 4934 || ((pixel_index2 >= 4994) && (pixel_index2 <= 4996)) || ((pixel_index2 >= 4998) && (pixel_index2 <= 5000)) || ((pixel_index2 >= 5021) && (pixel_index2 <= 5023)) || pixel_index2 == 5029 || ((pixel_index2 >= 5094) && (pixel_index2 <= 5096)) || ((pixel_index2 >= 5117) && (pixel_index2 <= 5118)) || ((pixel_index2 >= 5123) && (pixel_index2 <= 5124)) || ((pixel_index2 >= 5214) && (pixel_index2 <= 5218)) || ((pixel_index2 >= 5285) && (pixel_index2 <= 5286)) || ((pixel_index2 >= 5310) && (pixel_index2 <= 5313)) || ((pixel_index2 >= 5382) && (pixel_index2 <= 5383)) || ((pixel_index2 >= 5406) && (pixel_index2 <= 5407)) || ((pixel_index2 >= 5478) && (pixel_index2 <= 5479)) || pixel_index2 == 5503 || ((pixel_index2 >= 5573) && (pixel_index2 <= 5576)) || ((pixel_index2 >= 5584) && (pixel_index2 <= 5585)) || ((pixel_index2 >= 5591) && (pixel_index2 <= 5593)) || ((pixel_index2 >= 5598) && (pixel_index2 <= 5599)) || ((pixel_index2 >= 5671) && (pixel_index2 <= 5672)) || ((pixel_index2 >= 5680) && (pixel_index2 <= 5682)) || ((pixel_index2 >= 5687) && (pixel_index2 <= 5693)) || ((pixel_index2 >= 5777) && (pixel_index2 <= 5778)) || ((pixel_index2 >= 5785) && (pixel_index2 <= 5787)) || pixel_index2 == 5873 || pixel_index2 == 5969) oled_data2 = 16'b1010000000000000;
            else if (pixel_index2 == 5626 || pixel_index2 == 5630 || ((pixel_index2 >= 5634) && (pixel_index2 <= 5636)) || ((pixel_index2 >= 5638) && (pixel_index2 <= 5641)) || pixel_index2 == 5645 || pixel_index2 == 5649 || pixel_index2 == 5652 || ((pixel_index2 >= 5655) && (pixel_index2 <= 5656)) || ((pixel_index2 >= 5660) && (pixel_index2 <= 5662)) || pixel_index2 == 5729 || pixel_index2 == 5732 || pixel_index2 == 5737 || pixel_index2 == 5741 || pixel_index2 == 5746 || pixel_index2 == 5748 || pixel_index2 == 5750 || pixel_index2 == 5753 || pixel_index2 == 5755 || pixel_index2 == 5818 || pixel_index2 == 5822 || pixel_index2 == 5825 || pixel_index2 == 5828 || ((pixel_index2 >= 5831) && (pixel_index2 <= 5833)) || pixel_index2 == 5837 || ((pixel_index2 >= 5842) && (pixel_index2 <= 5844)) || pixel_index2 == 5846 || pixel_index2 == 5849 || ((pixel_index2 >= 5852) && (pixel_index2 <= 5853)) || pixel_index2 == 5914 || pixel_index2 == 5918 || pixel_index2 == 5921 || pixel_index2 == 5924 || pixel_index2 == 5929 || pixel_index2 == 5933 || pixel_index2 == 5937 || pixel_index2 == 5940 || pixel_index2 == 5942 || pixel_index2 == 5945 || pixel_index2 == 5950 || pixel_index2 == 6010 || pixel_index2 == 6014 || ((pixel_index2 >= 6018) && (pixel_index2 <= 6020)) || ((pixel_index2 >= 6022) && (pixel_index2 <= 6025)) || ((pixel_index2 >= 6027) && (pixel_index2 <= 6031)) || ((pixel_index2 >= 6034) && (pixel_index2 <= 6036)) || ((pixel_index2 >= 6039) && (pixel_index2 <= 6040)) || (pixel_index2 >= 6043) && (pixel_index2 <= 6045)) oled_data2 = 16'b0000000000010100;
            else oled_data2 = 0;
            end
            4: begin
            if (pixel_index2 == 163 || pixel_index2 == 356 || pixel_index2 == 643 || pixel_index2 == 740 || pixel_index2 == 836 || pixel_index2 == 932 || ((pixel_index2 >= 1221) && (pixel_index2 <= 1222)) || ((pixel_index2 >= 1318) && (pixel_index2 <= 1319)) || ((pixel_index2 >= 1414) && (pixel_index2 <= 1416)) || ((pixel_index2 >= 1510) && (pixel_index2 <= 1513)) || ((pixel_index2 >= 1607) && (pixel_index2 <= 1610)) || ((pixel_index2 >= 1703) && (pixel_index2 <= 1706)) || ((pixel_index2 >= 1800) && (pixel_index2 <= 1803)) || ((pixel_index2 >= 1896) && (pixel_index2 <= 1899)) || ((pixel_index2 >= 1992) && (pixel_index2 <= 1996)) || ((pixel_index2 >= 2089) && (pixel_index2 <= 2093)) || ((pixel_index2 >= 2185) && (pixel_index2 <= 2189)) || ((pixel_index2 >= 2281) && (pixel_index2 <= 2285)) || ((pixel_index2 >= 2378) && (pixel_index2 <= 2379)) || (pixel_index2 >= 2474) && (pixel_index2 <= 2475)) oled_data2 = 16'b1111001010000000;
            else if (pixel_index2 == 168 || ((pixel_index2 >= 172) && (pixel_index2 <= 175)) || ((pixel_index2 >= 178) && (pixel_index2 <= 180)) || ((pixel_index2 >= 182) && (pixel_index2 <= 185)) || pixel_index2 == 187 || pixel_index2 == 190 || pixel_index2 == 264 || pixel_index2 == 271 || pixel_index2 == 273 || pixel_index2 == 281 || pixel_index2 == 284 || pixel_index2 == 286 || pixel_index2 == 360 || ((pixel_index2 >= 365) && (pixel_index2 <= 367)) || ((pixel_index2 >= 370) && (pixel_index2 <= 371)) || ((pixel_index2 >= 375) && (pixel_index2 <= 377)) || ((pixel_index2 >= 380) && (pixel_index2 <= 382)) || pixel_index2 == 456 || pixel_index2 == 463 || pixel_index2 == 468 || pixel_index2 == 473 || pixel_index2 == 475 || pixel_index2 == 478 || ((pixel_index2 >= 550) && (pixel_index2 <= 554)) || ((pixel_index2 >= 556) && (pixel_index2 <= 559)) || ((pixel_index2 >= 561) && (pixel_index2 <= 563)) || ((pixel_index2 >= 566) && (pixel_index2 <= 569)) || ((pixel_index2 >= 572) && (pixel_index2 <= 574)) || ((pixel_index2 >= 744) && (pixel_index2 <= 746)) || ((pixel_index2 >= 749) && (pixel_index2 <= 751)) || ((pixel_index2 >= 753) && (pixel_index2 <= 756)) || pixel_index2 == 758 || pixel_index2 == 761 || pixel_index2 == 766 || pixel_index2 == 839 || pixel_index2 == 844 || pixel_index2 == 852 || pixel_index2 == 855 || pixel_index2 == 857 || pixel_index2 == 862 || ((pixel_index2 >= 936) && (pixel_index2 <= 937)) || ((pixel_index2 >= 941) && (pixel_index2 <= 942)) || ((pixel_index2 >= 946) && (pixel_index2 <= 948)) || ((pixel_index2 >= 951) && (pixel_index2 <= 953)) || ((pixel_index2 >= 956) && (pixel_index2 <= 958)) || pixel_index2 == 1034 || pixel_index2 == 1039 || pixel_index2 == 1044 || pixel_index2 == 1046 || pixel_index2 == 1049 || pixel_index2 == 1051 || pixel_index2 == 1054 || ((pixel_index2 >= 1127) && (pixel_index2 <= 1129)) || ((pixel_index2 >= 1132) && (pixel_index2 <= 1134)) || ((pixel_index2 >= 1137) && (pixel_index2 <= 1140)) || ((pixel_index2 >= 1143) && (pixel_index2 <= 1145)) || (pixel_index2 >= 1148) && (pixel_index2 <= 1150)) oled_data2 = 16'b1111010100000000;
            else if (((pixel_index2 >= 2380) && (pixel_index2 <= 2383)) || ((pixel_index2 >= 2476) && (pixel_index2 <= 2479)) || ((pixel_index2 >= 2572) && (pixel_index2 <= 2575)) || ((pixel_index2 >= 2668) && (pixel_index2 <= 2671)) || pixel_index2 == 3677 || pixel_index2 == 3760 || pixel_index2 == 3766 || pixel_index2 == 3942 || pixel_index2 == 3970 || pixel_index2 == 4321 || pixel_index2 == 4935 || pixel_index2 == 4993 || pixel_index2 == 5572 || pixel_index2 == 6065) oled_data2 = 16'b1111011110011110;
            else if (pixel_index2 == 3773 || ((pixel_index2 >= 3856) && (pixel_index2 <= 3857)) || pixel_index2 == 3862 || pixel_index2 == 3869 || pixel_index2 == 4038 || ((pixel_index2 >= 4065) && (pixel_index2 <= 4066)) || pixel_index2 == 4134 || pixel_index2 == 4161 || pixel_index2 == 4322 || pixel_index2 == 4934 || ((pixel_index2 >= 4994) && (pixel_index2 <= 4995)) || ((pixel_index2 >= 5029) && (pixel_index2 <= 5030)) || pixel_index2 == 5573 || pixel_index2 == 5873 || pixel_index2 == 5969) oled_data2 = 16'b1010000000000000;
            else if (pixel_index2 == 5626 || pixel_index2 == 5630 || ((pixel_index2 >= 5634) && (pixel_index2 <= 5636)) || ((pixel_index2 >= 5638) && (pixel_index2 <= 5641)) || pixel_index2 == 5645 || pixel_index2 == 5649 || pixel_index2 == 5652 || ((pixel_index2 >= 5655) && (pixel_index2 <= 5656)) || ((pixel_index2 >= 5660) && (pixel_index2 <= 5662)) || pixel_index2 == 5729 || pixel_index2 == 5732 || pixel_index2 == 5737 || pixel_index2 == 5741 || pixel_index2 == 5746 || pixel_index2 == 5748 || pixel_index2 == 5750 || pixel_index2 == 5753 || pixel_index2 == 5755 || pixel_index2 == 5818 || pixel_index2 == 5822 || pixel_index2 == 5825 || pixel_index2 == 5828 || ((pixel_index2 >= 5831) && (pixel_index2 <= 5833)) || pixel_index2 == 5837 || ((pixel_index2 >= 5842) && (pixel_index2 <= 5844)) || pixel_index2 == 5846 || pixel_index2 == 5849 || ((pixel_index2 >= 5852) && (pixel_index2 <= 5853)) || pixel_index2 == 5914 || pixel_index2 == 5918 || pixel_index2 == 5921 || pixel_index2 == 5924 || pixel_index2 == 5929 || pixel_index2 == 5933 || pixel_index2 == 5937 || pixel_index2 == 5940 || pixel_index2 == 5942 || pixel_index2 == 5945 || pixel_index2 == 5950 || pixel_index2 == 6010 || pixel_index2 == 6014 || ((pixel_index2 >= 6018) && (pixel_index2 <= 6020)) || ((pixel_index2 >= 6022) && (pixel_index2 <= 6025)) || ((pixel_index2 >= 6027) && (pixel_index2 <= 6031)) || ((pixel_index2 >= 6034) && (pixel_index2 <= 6036)) || ((pixel_index2 >= 6039) && (pixel_index2 <= 6040)) || (pixel_index2 >= 6043) && (pixel_index2 <= 6045)) oled_data2 = 16'b0000010100000000;
            else oled_data2 = 0;
            end
            5: begin
            if (((pixel_index2 >= 54) && (pixel_index2 <= 57)) || ((pixel_index2 >= 150) && (pixel_index2 <= 153)) || ((pixel_index2 >= 246) && (pixel_index2 <= 249)) || ((pixel_index2 >= 342) && (pixel_index2 <= 345)) || pixel_index2 == 3639 || ((pixel_index2 >= 3733) && (pixel_index2 <= 3736)) || ((pixel_index2 >= 3829) && (pixel_index2 <= 3832)) || ((pixel_index2 >= 3925) && (pixel_index2 <= 3928)) || (pixel_index2 >= 4021) && (pixel_index2 <= 4023)) oled_data2 = 16'b1111011110011110;
            else if (pixel_index2 == 168 || ((pixel_index2 >= 172) && (pixel_index2 <= 175)) || ((pixel_index2 >= 178) && (pixel_index2 <= 180)) || ((pixel_index2 >= 182) && (pixel_index2 <= 185)) || pixel_index2 == 187 || pixel_index2 == 190 || pixel_index2 == 264 || pixel_index2 == 271 || pixel_index2 == 273 || pixel_index2 == 281 || pixel_index2 == 284 || pixel_index2 == 286 || pixel_index2 == 360 || ((pixel_index2 >= 365) && (pixel_index2 <= 367)) || ((pixel_index2 >= 370) && (pixel_index2 <= 371)) || ((pixel_index2 >= 375) && (pixel_index2 <= 377)) || ((pixel_index2 >= 380) && (pixel_index2 <= 382)) || pixel_index2 == 456 || pixel_index2 == 463 || pixel_index2 == 468 || pixel_index2 == 473 || pixel_index2 == 475 || pixel_index2 == 478 || ((pixel_index2 >= 550) && (pixel_index2 <= 554)) || ((pixel_index2 >= 556) && (pixel_index2 <= 559)) || ((pixel_index2 >= 561) && (pixel_index2 <= 563)) || ((pixel_index2 >= 566) && (pixel_index2 <= 569)) || ((pixel_index2 >= 572) && (pixel_index2 <= 574)) || ((pixel_index2 >= 744) && (pixel_index2 <= 746)) || ((pixel_index2 >= 749) && (pixel_index2 <= 751)) || ((pixel_index2 >= 753) && (pixel_index2 <= 756)) || pixel_index2 == 758 || pixel_index2 == 761 || pixel_index2 == 766 || pixel_index2 == 839 || pixel_index2 == 844 || pixel_index2 == 852 || pixel_index2 == 855 || pixel_index2 == 857 || pixel_index2 == 862 || ((pixel_index2 >= 936) && (pixel_index2 <= 937)) || ((pixel_index2 >= 941) && (pixel_index2 <= 942)) || ((pixel_index2 >= 946) && (pixel_index2 <= 948)) || ((pixel_index2 >= 951) && (pixel_index2 <= 953)) || ((pixel_index2 >= 956) && (pixel_index2 <= 958)) || pixel_index2 == 1034 || pixel_index2 == 1039 || pixel_index2 == 1044 || pixel_index2 == 1046 || pixel_index2 == 1049 || pixel_index2 == 1051 || pixel_index2 == 1054 || ((pixel_index2 >= 1127) && (pixel_index2 <= 1129)) || ((pixel_index2 >= 1132) && (pixel_index2 <= 1134)) || ((pixel_index2 >= 1137) && (pixel_index2 <= 1140)) || ((pixel_index2 >= 1143) && (pixel_index2 <= 1145)) || (pixel_index2 >= 1148) && (pixel_index2 <= 1150)) oled_data2 = 16'b1111000000001010;
            else if (pixel_index2 == 1511 || pixel_index2 == 1704 || pixel_index2 == 1800 || pixel_index2 == 1900 || pixel_index2 == 1996 || ((pixel_index2 >= 2187) && (pixel_index2 <= 2188)) || ((pixel_index2 >= 2283) && (pixel_index2 <= 2286)) || ((pixel_index2 >= 2379) && (pixel_index2 <= 2382)) || ((pixel_index2 >= 2475) && (pixel_index2 <= 2478)) || ((pixel_index2 >= 2572) && (pixel_index2 <= 2575)) || ((pixel_index2 >= 2669) && (pixel_index2 <= 2672)) || ((pixel_index2 >= 2765) && (pixel_index2 <= 2769)) || ((pixel_index2 >= 2862) && (pixel_index2 <= 2866)) || ((pixel_index2 >= 2958) && (pixel_index2 <= 2962)) || ((pixel_index2 >= 3055) && (pixel_index2 <= 3059)) || ((pixel_index2 >= 3152) && (pixel_index2 <= 3155)) || ((pixel_index2 >= 3248) && (pixel_index2 <= 3252)) || ((pixel_index2 >= 3344) && (pixel_index2 <= 3349)) || ((pixel_index2 >= 3441) && (pixel_index2 <= 3446)) || ((pixel_index2 >= 3538) && (pixel_index2 <= 3542)) || ((pixel_index2 >= 3634) && (pixel_index2 <= 3637)) || ((pixel_index2 >= 3730) && (pixel_index2 <= 3732)) || (pixel_index2 >= 3827) && (pixel_index2 <= 3828)) oled_data2 = 16'b1111001010000000;
            else if (pixel_index2 == 5626 || pixel_index2 == 5630 || ((pixel_index2 >= 5634) && (pixel_index2 <= 5636)) || ((pixel_index2 >= 5638) && (pixel_index2 <= 5641)) || pixel_index2 == 5645 || pixel_index2 == 5649 || pixel_index2 == 5652 || ((pixel_index2 >= 5655) && (pixel_index2 <= 5656)) || ((pixel_index2 >= 5660) && (pixel_index2 <= 5662)) || pixel_index2 == 5729 || pixel_index2 == 5732 || pixel_index2 == 5737 || pixel_index2 == 5741 || pixel_index2 == 5746 || pixel_index2 == 5748 || pixel_index2 == 5750 || pixel_index2 == 5753 || pixel_index2 == 5755 || pixel_index2 == 5818 || pixel_index2 == 5822 || pixel_index2 == 5825 || pixel_index2 == 5828 || ((pixel_index2 >= 5831) && (pixel_index2 <= 5833)) || pixel_index2 == 5837 || ((pixel_index2 >= 5842) && (pixel_index2 <= 5844)) || pixel_index2 == 5846 || pixel_index2 == 5849 || ((pixel_index2 >= 5852) && (pixel_index2 <= 5853)) || pixel_index2 == 5914 || pixel_index2 == 5918 || pixel_index2 == 5921 || pixel_index2 == 5924 || pixel_index2 == 5929 || pixel_index2 == 5933 || pixel_index2 == 5937 || pixel_index2 == 5940 || pixel_index2 == 5942 || pixel_index2 == 5945 || pixel_index2 == 5950 || pixel_index2 == 6010 || pixel_index2 == 6014 || ((pixel_index2 >= 6018) && (pixel_index2 <= 6020)) || ((pixel_index2 >= 6022) && (pixel_index2 <= 6025)) || ((pixel_index2 >= 6027) && (pixel_index2 <= 6031)) || ((pixel_index2 >= 6034) && (pixel_index2 <= 6036)) || ((pixel_index2 >= 6039) && (pixel_index2 <= 6040)) || (pixel_index2 >= 6043) && (pixel_index2 <= 6045)) oled_data2 = 16'b1010000000000000;
            else oled_data2 = 0;
            end
            6: begin
            if (pixel_index2 == 168 || ((pixel_index2 >= 172) && (pixel_index2 <= 175)) || ((pixel_index2 >= 178) && (pixel_index2 <= 180)) || ((pixel_index2 >= 182) && (pixel_index2 <= 185)) || pixel_index2 == 187 || pixel_index2 == 190 || pixel_index2 == 264 || pixel_index2 == 271 || pixel_index2 == 273 || pixel_index2 == 281 || pixel_index2 == 284 || pixel_index2 == 286 || pixel_index2 == 360 || ((pixel_index2 >= 365) && (pixel_index2 <= 367)) || ((pixel_index2 >= 370) && (pixel_index2 <= 371)) || ((pixel_index2 >= 375) && (pixel_index2 <= 377)) || ((pixel_index2 >= 380) && (pixel_index2 <= 382)) || pixel_index2 == 456 || pixel_index2 == 463 || pixel_index2 == 468 || pixel_index2 == 473 || pixel_index2 == 475 || pixel_index2 == 478 || ((pixel_index2 >= 550) && (pixel_index2 <= 554)) || ((pixel_index2 >= 556) && (pixel_index2 <= 559)) || ((pixel_index2 >= 561) && (pixel_index2 <= 563)) || ((pixel_index2 >= 566) && (pixel_index2 <= 569)) || ((pixel_index2 >= 572) && (pixel_index2 <= 574)) || ((pixel_index2 >= 744) && (pixel_index2 <= 746)) || ((pixel_index2 >= 749) && (pixel_index2 <= 751)) || ((pixel_index2 >= 753) && (pixel_index2 <= 756)) || pixel_index2 == 758 || pixel_index2 == 761 || pixel_index2 == 766 || pixel_index2 == 839 || pixel_index2 == 844 || pixel_index2 == 852 || pixel_index2 == 855 || pixel_index2 == 857 || pixel_index2 == 862 || ((pixel_index2 >= 936) && (pixel_index2 <= 937)) || ((pixel_index2 >= 941) && (pixel_index2 <= 942)) || ((pixel_index2 >= 946) && (pixel_index2 <= 948)) || ((pixel_index2 >= 951) && (pixel_index2 <= 953)) || ((pixel_index2 >= 956) && (pixel_index2 <= 958)) || pixel_index2 == 1034 || pixel_index2 == 1039 || pixel_index2 == 1044 || pixel_index2 == 1046 || pixel_index2 == 1049 || pixel_index2 == 1051 || pixel_index2 == 1054 || ((pixel_index2 >= 1127) && (pixel_index2 <= 1129)) || ((pixel_index2 >= 1132) && (pixel_index2 <= 1134)) || ((pixel_index2 >= 1137) && (pixel_index2 <= 1140)) || ((pixel_index2 >= 1143) && (pixel_index2 <= 1145)) || (pixel_index2 >= 1148) && (pixel_index2 <= 1150)) oled_data2 = 16'b0000011110011110;
            else if (((pixel_index2 >= 247) && (pixel_index2 <= 248)) || ((pixel_index2 >= 342) && (pixel_index2 <= 344)) || pixel_index2 == 347 || ((pixel_index2 >= 437) && (pixel_index2 <= 439)) || ((pixel_index2 >= 533) && (pixel_index2 <= 535)) || pixel_index2 == 538 || ((pixel_index2 >= 628) && (pixel_index2 <= 630)) || pixel_index2 == 634 || ((pixel_index2 >= 722) && (pixel_index2 <= 725)) || ((pixel_index2 >= 817) && (pixel_index2 <= 821)) || ((pixel_index2 >= 912) && (pixel_index2 <= 915)) || ((pixel_index2 >= 1005) && (pixel_index2 <= 1011)) || ((pixel_index2 >= 1099) && (pixel_index2 <= 1106)) || ((pixel_index2 >= 1195) && (pixel_index2 <= 1201)) || ((pixel_index2 >= 1293) && (pixel_index2 <= 1295)) || (pixel_index2 >= 1389) && (pixel_index2 <= 1390)) oled_data2 = 16'b1111001010000000;
            else if (((pixel_index2 >= 1289) && (pixel_index2 <= 1292)) || ((pixel_index2 >= 1385) && (pixel_index2 <= 1388)) || ((pixel_index2 >= 1481) && (pixel_index2 <= 1484)) || ((pixel_index2 >= 1577) && (pixel_index2 <= 1580)) || ((pixel_index2 >= 2195) && (pixel_index2 <= 2196)) || ((pixel_index2 >= 2202) && (pixel_index2 <= 2203)) || ((pixel_index2 >= 2291) && (pixel_index2 <= 2292)) || ((pixel_index2 >= 2298) && (pixel_index2 <= 2299)) || ((pixel_index2 >= 2376) && (pixel_index2 <= 2377)) || ((pixel_index2 >= 2472) && (pixel_index2 <= 2473)) || ((pixel_index2 >= 2947) && (pixel_index2 <= 2948)) || ((pixel_index2 >= 3043) && (pixel_index2 <= 3044)) || pixel_index2 == 3734 || ((pixel_index2 >= 3811) && (pixel_index2 <= 3812)) || ((pixel_index2 >= 3829) && (pixel_index2 <= 3830)) || ((pixel_index2 >= 3907) && (pixel_index2 <= 3908)) || ((pixel_index2 >= 3924) && (pixel_index2 <= 3928)) || ((pixel_index2 >= 4019) && (pixel_index2 <= 4023)) || pixel_index2 == 4117 || ((pixel_index2 >= 4119) && (pixel_index2 <= 4120)) || ((pixel_index2 >= 4678) && (pixel_index2 <= 4679)) || ((pixel_index2 >= 4774) && (pixel_index2 <= 4775)) || ((pixel_index2 >= 5365) && (pixel_index2 <= 5366)) || (pixel_index2 >= 5461) && (pixel_index2 <= 5462)) oled_data2 = 16'b1111011110011110;
            else if (((pixel_index2 >= 2388) && (pixel_index2 <= 2389)) || pixel_index2 == 2394 || ((pixel_index2 >= 2484) && (pixel_index2 <= 2485)) || pixel_index2 == 2490 || ((pixel_index2 >= 2568) && (pixel_index2 <= 2569)) || ((pixel_index2 >= 2580) && (pixel_index2 <= 2581)) || pixel_index2 == 2586 || ((pixel_index2 >= 2664) && (pixel_index2 <= 2665)) || pixel_index2 == 2671 || pixel_index2 == 2677 || pixel_index2 == 2682 || pixel_index2 == 2761 || pixel_index2 == 2767 || pixel_index2 == 2773 || ((pixel_index2 >= 2777) && (pixel_index2 <= 2778)) || pixel_index2 == 2783 || pixel_index2 == 2855 || ((pixel_index2 >= 2857) && (pixel_index2 <= 2858)) || ((pixel_index2 >= 2863) && (pixel_index2 <= 2864)) || pixel_index2 == 2873 || pixel_index2 == 2879 || pixel_index2 == 2952 || ((pixel_index2 >= 2954) && (pixel_index2 <= 2957)) || pixel_index2 == 2960 || pixel_index2 == 2968 || pixel_index2 == 2974 || pixel_index2 == 3045 || pixel_index2 == 3048 || ((pixel_index2 >= 3051) && (pixel_index2 <= 3059)) || pixel_index2 == 3064 || ((pixel_index2 >= 3068) && (pixel_index2 <= 3069)) || pixel_index2 == 3142 || ((pixel_index2 >= 3147) && (pixel_index2 <= 3148)) || ((pixel_index2 >= 3153) && (pixel_index2 <= 3154)) || ((pixel_index2 >= 3159) && (pixel_index2 <= 3160)) || ((pixel_index2 >= 3162) && (pixel_index2 <= 3165)) || pixel_index2 == 3167 || pixel_index2 == 3239 || ((pixel_index2 >= 3245) && (pixel_index2 <= 3246)) || pixel_index2 == 3250 || pixel_index2 == 3259 || pixel_index2 == 3335 || pixel_index2 == 3346 || pixel_index2 == 3355 || pixel_index2 == 3431 || pixel_index2 == 3439 || pixel_index2 == 3442 || pixel_index2 == 3451 || ((pixel_index2 >= 3530) && (pixel_index2 <= 3533)) || pixel_index2 == 3535 || pixel_index2 == 3539 || pixel_index2 == 3547 || pixel_index2 == 3623 || pixel_index2 == 3631 || pixel_index2 == 3642 || ((pixel_index2 >= 3719) && (pixel_index2 <= 3720)) || pixel_index2 == 3738 || pixel_index2 == 3813 || ((pixel_index2 >= 3816) && (pixel_index2 <= 3817)) || ((pixel_index2 >= 3823) && (pixel_index2 <= 3824)) || ((pixel_index2 >= 3837) && (pixel_index2 <= 3839)) || ((pixel_index2 >= 3909) && (pixel_index2 <= 3911)) || ((pixel_index2 >= 3913) && (pixel_index2 <= 3914)) || ((pixel_index2 >= 3916) && (pixel_index2 <= 3917)) || pixel_index2 == 3920 || ((pixel_index2 >= 3933) && (pixel_index2 <= 3934)) || ((pixel_index2 >= 4028) && (pixel_index2 <= 4029)) || ((pixel_index2 >= 4200) && (pixel_index2 <= 4201)) || ((pixel_index2 >= 4296) && (pixel_index2 <= 4297)) || ((pixel_index2 >= 4302) && (pixel_index2 <= 4304)) || ((pixel_index2 >= 4392) && (pixel_index2 <= 4393)) || ((pixel_index2 >= 4398) && (pixel_index2 <= 4401)) || ((pixel_index2 >= 4489) && (pixel_index2 <= 4491)) || ((pixel_index2 >= 4500) && (pixel_index2 <= 4502)) || pixel_index2 == 4593 || pixel_index2 == 4595 || pixel_index2 == 4599 || ((pixel_index2 >= 4680) && (pixel_index2 <= 4681)) || pixel_index2 == 4689 || pixel_index2 == 4693 || pixel_index2 == 4696 || ((pixel_index2 >= 4698) && (pixel_index2 <= 4699)) || ((pixel_index2 >= 4792) && (pixel_index2 <= 4797)) || pixel_index2 == 4885 || ((pixel_index2 >= 4893) && (pixel_index2 <= 4895)) || pixel_index2 == 4981 || pixel_index2 == 5077 || pixel_index2 == 5173 || pixel_index2 == 5269 || pixel_index2 == 5626 || pixel_index2 == 5630 || ((pixel_index2 >= 5634) && (pixel_index2 <= 5636)) || ((pixel_index2 >= 5638) && (pixel_index2 <= 5641)) || pixel_index2 == 5645 || pixel_index2 == 5649 || pixel_index2 == 5652 || ((pixel_index2 >= 5655) && (pixel_index2 <= 5656)) || ((pixel_index2 >= 5660) && (pixel_index2 <= 5662)) || pixel_index2 == 5729 || pixel_index2 == 5732 || pixel_index2 == 5737 || pixel_index2 == 5741 || pixel_index2 == 5746 || pixel_index2 == 5748 || pixel_index2 == 5750 || pixel_index2 == 5753 || pixel_index2 == 5755 || pixel_index2 == 5818 || pixel_index2 == 5822 || pixel_index2 == 5825 || pixel_index2 == 5828 || ((pixel_index2 >= 5831) && (pixel_index2 <= 5833)) || pixel_index2 == 5837 || ((pixel_index2 >= 5842) && (pixel_index2 <= 5844)) || pixel_index2 == 5846 || pixel_index2 == 5849 || ((pixel_index2 >= 5852) && (pixel_index2 <= 5853)) || pixel_index2 == 5914 || pixel_index2 == 5918 || pixel_index2 == 5921 || pixel_index2 == 5924 || pixel_index2 == 5929 || pixel_index2 == 5933 || pixel_index2 == 5937 || pixel_index2 == 5940 || pixel_index2 == 5942 || pixel_index2 == 5945 || pixel_index2 == 5950 || pixel_index2 == 6010 || pixel_index2 == 6014 || ((pixel_index2 >= 6018) && (pixel_index2 <= 6020)) || ((pixel_index2 >= 6022) && (pixel_index2 <= 6025)) || ((pixel_index2 >= 6027) && (pixel_index2 <= 6031)) || ((pixel_index2 >= 6034) && (pixel_index2 <= 6036)) || ((pixel_index2 >= 6039) && (pixel_index2 <= 6040)) || (pixel_index2 >= 6043) && (pixel_index2 <= 6045)) oled_data2 = 16'b0000000000010100;
            else if (pixel_index2 == 2965 || pixel_index2 == 3061 || pixel_index2 == 3157 || pixel_index2 == 3247 || pixel_index2 == 3253 || pixel_index2 == 3258 || ((pixel_index2 >= 3343) && (pixel_index2 <= 3344)) || pixel_index2 == 3349 || pixel_index2 == 3354 || ((pixel_index2 >= 3440) && (pixel_index2 <= 3441)) || pixel_index2 == 3445 || pixel_index2 == 3450 || ((pixel_index2 >= 3537) && (pixel_index2 <= 3538)) || ((pixel_index2 >= 3540) && (pixel_index2 <= 3546)) || pixel_index2 == 3550 || ((pixel_index2 >= 3628) && (pixel_index2 <= 3630)) || ((pixel_index2 >= 3632) && (pixel_index2 <= 3641)) || ((pixel_index2 >= 3644) && (pixel_index2 <= 3646)) || ((pixel_index2 >= 3726) && (pixel_index2 <= 3733)) || ((pixel_index2 >= 3735) && (pixel_index2 <= 3737)) || ((pixel_index2 >= 3739) && (pixel_index2 <= 3741)) || ((pixel_index2 >= 3825) && (pixel_index2 <= 3828)) || ((pixel_index2 >= 3831) && (pixel_index2 <= 3836)) || ((pixel_index2 >= 3918) && (pixel_index2 <= 3919)) || ((pixel_index2 >= 3921) && (pixel_index2 <= 3923)) || ((pixel_index2 >= 3929) && (pixel_index2 <= 3932)) || ((pixel_index2 >= 4011) && (pixel_index2 <= 4018)) || ((pixel_index2 >= 4024) && (pixel_index2 <= 4027)) || ((pixel_index2 >= 4108) && (pixel_index2 <= 4116)) || pixel_index2 == 4118 || ((pixel_index2 >= 4121) && (pixel_index2 <= 4123)) || pixel_index2 == 4125 || ((pixel_index2 >= 4205) && (pixel_index2 <= 4221)) || ((pixel_index2 >= 4305) && (pixel_index2 <= 4314)) || ((pixel_index2 >= 4402) && (pixel_index2 <= 4410)) || ((pixel_index2 >= 4498) && (pixel_index2 <= 4499)) || ((pixel_index2 >= 4503) && (pixel_index2 <= 4508)) || pixel_index2 == 4594 || ((pixel_index2 >= 4600) && (pixel_index2 <= 4605)) || pixel_index2 == 4690 || pixel_index2 == 4697) oled_data2 = 16'b1010010100011110;
            else oled_data2 = 0;
            end
            7: begin
            if (pixel_index2 == 168 || ((pixel_index2 >= 172) && (pixel_index2 <= 175)) || ((pixel_index2 >= 178) && (pixel_index2 <= 180)) || ((pixel_index2 >= 182) && (pixel_index2 <= 185)) || pixel_index2 == 187 || pixel_index2 == 190 || pixel_index2 == 264 || pixel_index2 == 271 || pixel_index2 == 273 || pixel_index2 == 281 || pixel_index2 == 284 || pixel_index2 == 286 || pixel_index2 == 360 || ((pixel_index2 >= 365) && (pixel_index2 <= 367)) || ((pixel_index2 >= 370) && (pixel_index2 <= 371)) || ((pixel_index2 >= 375) && (pixel_index2 <= 377)) || ((pixel_index2 >= 380) && (pixel_index2 <= 382)) || pixel_index2 == 456 || pixel_index2 == 463 || pixel_index2 == 468 || pixel_index2 == 473 || pixel_index2 == 475 || pixel_index2 == 478 || ((pixel_index2 >= 550) && (pixel_index2 <= 554)) || ((pixel_index2 >= 556) && (pixel_index2 <= 559)) || ((pixel_index2 >= 561) && (pixel_index2 <= 563)) || ((pixel_index2 >= 566) && (pixel_index2 <= 569)) || ((pixel_index2 >= 572) && (pixel_index2 <= 574)) || ((pixel_index2 >= 744) && (pixel_index2 <= 746)) || ((pixel_index2 >= 749) && (pixel_index2 <= 751)) || ((pixel_index2 >= 753) && (pixel_index2 <= 756)) || pixel_index2 == 758 || pixel_index2 == 761 || pixel_index2 == 766 || pixel_index2 == 839 || pixel_index2 == 844 || pixel_index2 == 852 || pixel_index2 == 855 || pixel_index2 == 857 || pixel_index2 == 862 || ((pixel_index2 >= 936) && (pixel_index2 <= 937)) || ((pixel_index2 >= 941) && (pixel_index2 <= 942)) || ((pixel_index2 >= 946) && (pixel_index2 <= 948)) || ((pixel_index2 >= 951) && (pixel_index2 <= 953)) || ((pixel_index2 >= 956) && (pixel_index2 <= 958)) || pixel_index2 == 1034 || pixel_index2 == 1039 || pixel_index2 == 1044 || pixel_index2 == 1046 || pixel_index2 == 1049 || pixel_index2 == 1051 || pixel_index2 == 1054 || ((pixel_index2 >= 1127) && (pixel_index2 <= 1129)) || ((pixel_index2 >= 1132) && (pixel_index2 <= 1134)) || ((pixel_index2 >= 1137) && (pixel_index2 <= 1140)) || ((pixel_index2 >= 1143) && (pixel_index2 <= 1145)) || (pixel_index2 >= 1148) && (pixel_index2 <= 1150)) oled_data2 = 16'b1111010100000000;
            else if (((pixel_index2 >= 1007) && (pixel_index2 <= 1008)) || ((pixel_index2 >= 1100) && (pixel_index2 <= 1103)) || ((pixel_index2 >= 1196) && (pixel_index2 <= 1198)) || pixel_index2 == 1202 || ((pixel_index2 >= 1291) && (pixel_index2 <= 1294)) || ((pixel_index2 >= 1383) && (pixel_index2 <= 1389)) || pixel_index2 == 1393 || pixel_index2 == 1475 || ((pixel_index2 >= 1478) && (pixel_index2 <= 1483)) || pixel_index2 == 1488 || ((pixel_index2 >= 1569) && (pixel_index2 <= 1577)) || ((pixel_index2 >= 1664) && (pixel_index2 <= 1673)) || ((pixel_index2 >= 1762) && (pixel_index2 <= 1766)) || (pixel_index2 >= 1858) && (pixel_index2 <= 1860)) oled_data2 = 16'b1111001010000000;
            else if (pixel_index2 == 1663 || ((pixel_index2 >= 1758) && (pixel_index2 <= 1761)) || ((pixel_index2 >= 1854) && (pixel_index2 <= 1857)) || ((pixel_index2 >= 1950) && (pixel_index2 <= 1953)) || ((pixel_index2 >= 2046) && (pixel_index2 <= 2049)) || ((pixel_index2 >= 2195) && (pixel_index2 <= 2196)) || ((pixel_index2 >= 2202) && (pixel_index2 <= 2203)) || ((pixel_index2 >= 2291) && (pixel_index2 <= 2292)) || ((pixel_index2 >= 2298) && (pixel_index2 <= 2299)) || ((pixel_index2 >= 2376) && (pixel_index2 <= 2377)) || ((pixel_index2 >= 2472) && (pixel_index2 <= 2473)) || ((pixel_index2 >= 2947) && (pixel_index2 <= 2948)) || ((pixel_index2 >= 3043) && (pixel_index2 <= 3044)) || ((pixel_index2 >= 3811) && (pixel_index2 <= 3812)) || ((pixel_index2 >= 3907) && (pixel_index2 <= 3908)) || ((pixel_index2 >= 4678) && (pixel_index2 <= 4679)) || ((pixel_index2 >= 4774) && (pixel_index2 <= 4775)) || ((pixel_index2 >= 5365) && (pixel_index2 <= 5366)) || (pixel_index2 >= 5461) && (pixel_index2 <= 5462)) oled_data2 = 16'b1111011110011110;
            else if (((pixel_index2 >= 2388) && (pixel_index2 <= 2389)) || pixel_index2 == 2394 || ((pixel_index2 >= 2484) && (pixel_index2 <= 2485)) || pixel_index2 == 2490 || ((pixel_index2 >= 2568) && (pixel_index2 <= 2569)) || ((pixel_index2 >= 2580) && (pixel_index2 <= 2581)) || pixel_index2 == 2586 || ((pixel_index2 >= 2664) && (pixel_index2 <= 2665)) || pixel_index2 == 2671 || pixel_index2 == 2677 || pixel_index2 == 2682 || pixel_index2 == 2761 || pixel_index2 == 2767 || ((pixel_index2 >= 2772) && (pixel_index2 <= 2773)) || ((pixel_index2 >= 2777) && (pixel_index2 <= 2778)) || pixel_index2 == 2783 || pixel_index2 == 2855 || ((pixel_index2 >= 2857) && (pixel_index2 <= 2858)) || ((pixel_index2 >= 2863) && (pixel_index2 <= 2864)) || ((pixel_index2 >= 2868) && (pixel_index2 <= 2869)) || ((pixel_index2 >= 2872) && (pixel_index2 <= 2874)) || pixel_index2 == 2879 || ((pixel_index2 >= 2952) && (pixel_index2 <= 2955)) || pixel_index2 == 2960 || ((pixel_index2 >= 2968) && (pixel_index2 <= 2969)) || pixel_index2 == 2974 || pixel_index2 == 3045 || ((pixel_index2 >= 3048) && (pixel_index2 <= 3051)) || ((pixel_index2 >= 3055) && (pixel_index2 <= 3057)) || ((pixel_index2 >= 3068) && (pixel_index2 <= 3070)) || pixel_index2 == 3142 || ((pixel_index2 >= 3146) && (pixel_index2 <= 3147)) || ((pixel_index2 >= 3151) && (pixel_index2 <= 3153)) || ((pixel_index2 >= 3164) && (pixel_index2 <= 3167)) || pixel_index2 == 3239 || ((pixel_index2 >= 3247) && (pixel_index2 <= 3248)) || ((pixel_index2 >= 3261) && (pixel_index2 <= 3262)) || pixel_index2 == 3335 || pixel_index2 == 3431 || pixel_index2 == 3623 || ((pixel_index2 >= 3719) && (pixel_index2 <= 3720)) || pixel_index2 == 3813 || ((pixel_index2 >= 3816) && (pixel_index2 <= 3817)) || ((pixel_index2 >= 3909) && (pixel_index2 <= 3914)) || ((pixel_index2 >= 4008) && (pixel_index2 <= 4010)) || ((pixel_index2 >= 4105) && (pixel_index2 <= 4106)) || pixel_index2 == 4392 || ((pixel_index2 >= 4489) && (pixel_index2 <= 4493)) || ((pixel_index2 >= 4586) && (pixel_index2 <= 4589)) || ((pixel_index2 >= 4680) && (pixel_index2 <= 4685)) || ((pixel_index2 >= 4699) && (pixel_index2 <= 4700)) || ((pixel_index2 >= 4778) && (pixel_index2 <= 4779)) || ((pixel_index2 >= 4788) && (pixel_index2 <= 4790)) || ((pixel_index2 >= 4795) && (pixel_index2 <= 4797)) || ((pixel_index2 >= 4884) && (pixel_index2 <= 4886)) || ((pixel_index2 >= 4893) && (pixel_index2 <= 4895)) || pixel_index2 == 4981 || pixel_index2 == 5077 || pixel_index2 == 5173 || pixel_index2 == 5269) oled_data2 = 16'b0000000000010100;
            else if (pixel_index2 == 5626 || pixel_index2 == 5630 || ((pixel_index2 >= 5634) && (pixel_index2 <= 5636)) || ((pixel_index2 >= 5638) && (pixel_index2 <= 5641)) || pixel_index2 == 5645 || pixel_index2 == 5649 || pixel_index2 == 5652 || ((pixel_index2 >= 5655) && (pixel_index2 <= 5656)) || ((pixel_index2 >= 5660) && (pixel_index2 <= 5662)) || pixel_index2 == 5729 || pixel_index2 == 5732 || pixel_index2 == 5737 || pixel_index2 == 5741 || pixel_index2 == 5746 || pixel_index2 == 5748 || pixel_index2 == 5750 || pixel_index2 == 5753 || pixel_index2 == 5755 || pixel_index2 == 5818 || pixel_index2 == 5822 || pixel_index2 == 5825 || pixel_index2 == 5828 || ((pixel_index2 >= 5831) && (pixel_index2 <= 5833)) || pixel_index2 == 5837 || ((pixel_index2 >= 5842) && (pixel_index2 <= 5844)) || pixel_index2 == 5846 || pixel_index2 == 5849 || ((pixel_index2 >= 5852) && (pixel_index2 <= 5853)) || pixel_index2 == 5914 || pixel_index2 == 5918 || pixel_index2 == 5921 || pixel_index2 == 5924 || pixel_index2 == 5929 || pixel_index2 == 5933 || pixel_index2 == 5937 || pixel_index2 == 5940 || pixel_index2 == 5942 || pixel_index2 == 5945 || pixel_index2 == 5950 || pixel_index2 == 6010 || pixel_index2 == 6014 || ((pixel_index2 >= 6018) && (pixel_index2 <= 6020)) || ((pixel_index2 >= 6022) && (pixel_index2 <= 6025)) || ((pixel_index2 >= 6027) && (pixel_index2 <= 6031)) || ((pixel_index2 >= 6034) && (pixel_index2 <= 6036)) || ((pixel_index2 >= 6039) && (pixel_index2 <= 6040)) || (pixel_index2 >= 6043) && (pixel_index2 <= 6045)) oled_data2 = 16'b0000010100000000;
            else oled_data2 = 0;
            end
            8: begin
            if (pixel_index2 == 168 || ((pixel_index2 >= 172) && (pixel_index2 <= 175)) || ((pixel_index2 >= 178) && (pixel_index2 <= 180)) || ((pixel_index2 >= 182) && (pixel_index2 <= 184)) || pixel_index2 == 187 || pixel_index2 == 264 || pixel_index2 == 271 || pixel_index2 == 273 || pixel_index2 == 284 || pixel_index2 == 360 || ((pixel_index2 >= 365) && (pixel_index2 <= 367)) || ((pixel_index2 >= 370) && (pixel_index2 <= 371)) || ((pixel_index2 >= 375) && (pixel_index2 <= 376)) || ((pixel_index2 >= 380) && (pixel_index2 <= 381)) || pixel_index2 == 456 || pixel_index2 == 463 || pixel_index2 == 468 || pixel_index2 == 475 || ((pixel_index2 >= 550) && (pixel_index2 <= 554)) || ((pixel_index2 >= 556) && (pixel_index2 <= 559)) || ((pixel_index2 >= 561) && (pixel_index2 <= 563)) || ((pixel_index2 >= 566) && (pixel_index2 <= 568)) || ((pixel_index2 >= 572) && (pixel_index2 <= 573)) || ((pixel_index2 >= 744) && (pixel_index2 <= 746)) || ((pixel_index2 >= 749) && (pixel_index2 <= 751)) || ((pixel_index2 >= 753) && (pixel_index2 <= 756)) || pixel_index2 == 758 || pixel_index2 == 839 || pixel_index2 == 844 || pixel_index2 == 852 || pixel_index2 == 855 || ((pixel_index2 >= 936) && (pixel_index2 <= 937)) || ((pixel_index2 >= 941) && (pixel_index2 <= 942)) || ((pixel_index2 >= 946) && (pixel_index2 <= 948)) || ((pixel_index2 >= 951) && (pixel_index2 <= 952)) || ((pixel_index2 >= 956) && (pixel_index2 <= 957)) || pixel_index2 == 1034 || pixel_index2 == 1039 || pixel_index2 == 1044 || pixel_index2 == 1046 || pixel_index2 == 1051 || ((pixel_index2 >= 1127) && (pixel_index2 <= 1129)) || ((pixel_index2 >= 1132) && (pixel_index2 <= 1134)) || ((pixel_index2 >= 1137) && (pixel_index2 <= 1140)) || ((pixel_index2 >= 1143) && (pixel_index2 <= 1144)) || (pixel_index2 >= 1148) && (pixel_index2 <= 1149)) oled_data2 = 16'b1111000000001010;
            else if (pixel_index2 == 185 || pixel_index2 == 190 || pixel_index2 == 281 || pixel_index2 == 286 || pixel_index2 == 377 || pixel_index2 == 382 || pixel_index2 == 473 || pixel_index2 == 478 || pixel_index2 == 569 || pixel_index2 == 574 || pixel_index2 == 761 || pixel_index2 == 766 || pixel_index2 == 857 || pixel_index2 == 862 || pixel_index2 == 953 || pixel_index2 == 958 || pixel_index2 == 1049 || pixel_index2 == 1054 || pixel_index2 == 1145 || pixel_index2 == 1150) oled_data2 = 16'b1010000000001010;
            else if (pixel_index2 == 186 || pixel_index2 == 474 || pixel_index2 == 1050 || pixel_index2 == 5754 || pixel_index2 == 6042) oled_data2 = 16'b0101000000000000;
            else if (((pixel_index2 >= 986) && (pixel_index2 <= 987)) || ((pixel_index2 >= 992) && (pixel_index2 <= 993)) || ((pixel_index2 >= 998) && (pixel_index2 <= 999)) || ((pixel_index2 >= 1082) && (pixel_index2 <= 1083)) || ((pixel_index2 >= 1088) && (pixel_index2 <= 1089)) || ((pixel_index2 >= 1094) && (pixel_index2 <= 1095)) || ((pixel_index2 >= 1194) && (pixel_index2 <= 1195)) || ((pixel_index2 >= 1267) && (pixel_index2 <= 1268)) || ((pixel_index2 >= 1290) && (pixel_index2 <= 1291)) || ((pixel_index2 >= 1363) && (pixel_index2 <= 1364)) || ((pixel_index2 >= 1465) && (pixel_index2 <= 1466)) || ((pixel_index2 >= 1471) && (pixel_index2 <= 1472)) || pixel_index2 == 1475 || ((pixel_index2 >= 1561) && (pixel_index2 <= 1563)) || ((pixel_index2 >= 1566) && (pixel_index2 <= 1568)) || ((pixel_index2 >= 1570) && (pixel_index2 <= 1571)) || ((pixel_index2 >= 1574) && (pixel_index2 <= 1575)) || pixel_index2 == 1655 || ((pixel_index2 >= 1658) && (pixel_index2 <= 1666)) || ((pixel_index2 >= 1669) && (pixel_index2 <= 1670)) || ((pixel_index2 >= 1742) && (pixel_index2 <= 1743)) || ((pixel_index2 >= 1751) && (pixel_index2 <= 1753)) || ((pixel_index2 >= 1755) && (pixel_index2 <= 1765)) || ((pixel_index2 >= 1838) && (pixel_index2 <= 1839)) || ((pixel_index2 >= 1848) && (pixel_index2 <= 1860)) || ((pixel_index2 >= 1868) && (pixel_index2 <= 1869)) || ((pixel_index2 >= 1945) && (pixel_index2 <= 1955)) || ((pixel_index2 >= 1964) && (pixel_index2 <= 1965)) || ((pixel_index2 >= 2043) && (pixel_index2 <= 2053)) || ((pixel_index2 >= 2138) && (pixel_index2 <= 2150)) || ((pixel_index2 >= 2231) && (pixel_index2 <= 2241)) || pixel_index2 == 2292 || ((pixel_index2 >= 2323) && (pixel_index2 <= 2324)) || ((pixel_index2 >= 2333) && (pixel_index2 <= 2335)) || ((pixel_index2 >= 2337) && (pixel_index2 <= 2338)) || ((pixel_index2 >= 2346) && (pixel_index2 <= 2347)) || ((pixel_index2 >= 2419) && (pixel_index2 <= 2420)) || pixel_index2 == 2429 || ((pixel_index2 >= 2442) && (pixel_index2 <= 2443)) || pixel_index2 == 2472 || ((pixel_index2 >= 2630) && (pixel_index2 <= 2631)) || ((pixel_index2 >= 2726) && (pixel_index2 <= 2727)) || ((pixel_index2 >= 2812) && (pixel_index2 <= 2813)) || ((pixel_index2 >= 2818) && (pixel_index2 <= 2819)) || ((pixel_index2 >= 2908) && (pixel_index2 <= 2909)) || ((pixel_index2 >= 2914) && (pixel_index2 <= 2915)) || pixel_index2 == 3044 || pixel_index2 == 3812 || pixel_index2 == 4679 || pixel_index2 == 5365) oled_data2 = 16'b1111011110011110;
            else if (pixel_index2 == 2298) oled_data2 = 16'b0101001010001010;
            else if (pixel_index2 == 2388 || pixel_index2 == 2485 || pixel_index2 == 2568 || pixel_index2 == 2664 || pixel_index2 == 2671 || pixel_index2 == 2772 || pixel_index2 == 2855 || pixel_index2 == 2864 || pixel_index2 == 2868 || pixel_index2 == 2872 || pixel_index2 == 2952 || pixel_index2 == 2955 || pixel_index2 == 3045 || pixel_index2 == 3048 || pixel_index2 == 3057 || pixel_index2 == 3068 || pixel_index2 == 3146 || pixel_index2 == 3153 || pixel_index2 == 3166 || pixel_index2 == 3248 || pixel_index2 == 3261 || pixel_index2 == 3335 || pixel_index2 == 3431 || pixel_index2 == 3623 || pixel_index2 == 3719 || pixel_index2 == 3813 || ((pixel_index2 >= 3909) && (pixel_index2 <= 3910)) || ((pixel_index2 >= 3913) && (pixel_index2 <= 3914)) || pixel_index2 == 4392 || ((pixel_index2 >= 4489) && (pixel_index2 <= 4492)) || pixel_index2 == 4680 || pixel_index2 == 4699 || pixel_index2 == 4778 || pixel_index2 == 4894 || pixel_index2 == 4981 || pixel_index2 == 5173 || pixel_index2 == 5269) oled_data2 = 16'b0000000000010100;
            else if (pixel_index2 == 2394 || pixel_index2 == 2490 || pixel_index2 == 2586 || pixel_index2 == 2777 || pixel_index2 == 2783 || pixel_index2 == 2873 || pixel_index2 == 2879 || pixel_index2 == 2968 || pixel_index2 == 3167 || pixel_index2 == 3262 || pixel_index2 == 4698 || pixel_index2 == 4895) oled_data2 = 16'b0000000000001010;
            else if (pixel_index2 == 5626 || pixel_index2 == 5630 || ((pixel_index2 >= 5634) && (pixel_index2 <= 5636)) || ((pixel_index2 >= 5638) && (pixel_index2 <= 5641)) || pixel_index2 == 5645 || pixel_index2 == 5649 || pixel_index2 == 5652 || ((pixel_index2 >= 5655) && (pixel_index2 <= 5656)) || ((pixel_index2 >= 5660) && (pixel_index2 <= 5662)) || pixel_index2 == 5729 || pixel_index2 == 5732 || pixel_index2 == 5737 || pixel_index2 == 5741 || pixel_index2 == 5746 || pixel_index2 == 5748 || pixel_index2 == 5750 || pixel_index2 == 5753 || pixel_index2 == 5755 || pixel_index2 == 5818 || pixel_index2 == 5822 || pixel_index2 == 5825 || pixel_index2 == 5828 || ((pixel_index2 >= 5831) && (pixel_index2 <= 5833)) || pixel_index2 == 5837 || ((pixel_index2 >= 5842) && (pixel_index2 <= 5844)) || pixel_index2 == 5846 || pixel_index2 == 5849 || ((pixel_index2 >= 5852) && (pixel_index2 <= 5853)) || pixel_index2 == 5914 || pixel_index2 == 5918 || pixel_index2 == 5921 || pixel_index2 == 5924 || pixel_index2 == 5929 || pixel_index2 == 5933 || pixel_index2 == 5937 || pixel_index2 == 5940 || pixel_index2 == 5942 || pixel_index2 == 5945 || pixel_index2 == 5950 || pixel_index2 == 6010 || pixel_index2 == 6014 || ((pixel_index2 >= 6018) && (pixel_index2 <= 6020)) || ((pixel_index2 >= 6022) && (pixel_index2 <= 6025)) || ((pixel_index2 >= 6027) && (pixel_index2 <= 6031)) || ((pixel_index2 >= 6034) && (pixel_index2 <= 6036)) || ((pixel_index2 >= 6039) && (pixel_index2 <= 6040)) || (pixel_index2 >= 6043) && (pixel_index2 <= 6045)) oled_data2 = 16'b1010000000000000;
            else oled_data2 = 0;
            end
            9: begin
            if (((pixel_index2 >= 138) && (pixel_index2 <= 139)) || ((pixel_index2 >= 217) && (pixel_index2 <= 218)) || ((pixel_index2 >= 225) && (pixel_index2 <= 226)) || ((pixel_index2 >= 234) && (pixel_index2 <= 235)) || ((pixel_index2 >= 313) && (pixel_index2 <= 314)) || ((pixel_index2 >= 321) && (pixel_index2 <= 322)) || ((pixel_index2 >= 494) && (pixel_index2 <= 495)) || ((pixel_index2 >= 527) && (pixel_index2 <= 528)) || ((pixel_index2 >= 590) && (pixel_index2 <= 591)) || ((pixel_index2 >= 623) && (pixel_index2 <= 624)) || ((pixel_index2 >= 1065) && (pixel_index2 <= 1066)) || ((pixel_index2 >= 1161) && (pixel_index2 <= 1162)) || ((pixel_index2 >= 1569) && (pixel_index2 <= 1570)) || ((pixel_index2 >= 1665) && (pixel_index2 <= 1666)) || ((pixel_index2 >= 1760) && (pixel_index2 <= 1762)) || ((pixel_index2 >= 1853) && (pixel_index2 <= 1859)) || ((pixel_index2 >= 1877) && (pixel_index2 <= 1878)) || ((pixel_index2 >= 1948) && (pixel_index2 <= 1958)) || ((pixel_index2 >= 1973) && (pixel_index2 <= 1974)) || ((pixel_index2 >= 2025) && (pixel_index2 <= 2026)) || ((pixel_index2 >= 2042) && (pixel_index2 <= 2055)) || ((pixel_index2 >= 2121) && (pixel_index2 <= 2122)) || ((pixel_index2 >= 2138) && (pixel_index2 <= 2150)) || ((pixel_index2 >= 2235) && (pixel_index2 <= 2244)) || ((pixel_index2 >= 2330) && (pixel_index2 <= 2338)) || ((pixel_index2 >= 2340) && (pixel_index2 <= 2341)) || ((pixel_index2 >= 2427) && (pixel_index2 <= 2433)) || ((pixel_index2 >= 2523) && (pixel_index2 <= 2528)) || ((pixel_index2 >= 2621) && (pixel_index2 <= 2624)) || pixel_index2 == 2719 || ((pixel_index2 >= 2833) && (pixel_index2 <= 2834)) || ((pixel_index2 >= 2929) && (pixel_index2 <= 2930)) || ((pixel_index2 >= 3084) && (pixel_index2 <= 3085)) || ((pixel_index2 >= 3180) && (pixel_index2 <= 3181)) || ((pixel_index2 >= 3593) && (pixel_index2 <= 3594)) || ((pixel_index2 >= 3676) && (pixel_index2 <= 3677)) || ((pixel_index2 >= 3689) && (pixel_index2 <= 3690)) || (pixel_index2 >= 3772) && (pixel_index2 <= 3773)) oled_data2 = 16'b1111011110011110;
            else if (pixel_index2 == 168 || ((pixel_index2 >= 172) && (pixel_index2 <= 175)) || ((pixel_index2 >= 178) && (pixel_index2 <= 180)) || ((pixel_index2 >= 182) && (pixel_index2 <= 185)) || pixel_index2 == 187 || pixel_index2 == 190 || pixel_index2 == 264 || pixel_index2 == 271 || pixel_index2 == 273 || pixel_index2 == 281 || pixel_index2 == 284 || pixel_index2 == 286 || pixel_index2 == 360 || ((pixel_index2 >= 365) && (pixel_index2 <= 367)) || ((pixel_index2 >= 370) && (pixel_index2 <= 371)) || ((pixel_index2 >= 375) && (pixel_index2 <= 377)) || ((pixel_index2 >= 380) && (pixel_index2 <= 382)) || pixel_index2 == 456 || pixel_index2 == 463 || pixel_index2 == 468 || pixel_index2 == 473 || pixel_index2 == 475 || pixel_index2 == 478 || ((pixel_index2 >= 550) && (pixel_index2 <= 554)) || ((pixel_index2 >= 556) && (pixel_index2 <= 559)) || ((pixel_index2 >= 561) && (pixel_index2 <= 563)) || ((pixel_index2 >= 566) && (pixel_index2 <= 569)) || ((pixel_index2 >= 572) && (pixel_index2 <= 574)) || ((pixel_index2 >= 744) && (pixel_index2 <= 746)) || ((pixel_index2 >= 749) && (pixel_index2 <= 751)) || ((pixel_index2 >= 753) && (pixel_index2 <= 756)) || pixel_index2 == 758 || pixel_index2 == 761 || pixel_index2 == 766 || pixel_index2 == 839 || pixel_index2 == 844 || pixel_index2 == 852 || pixel_index2 == 855 || pixel_index2 == 857 || pixel_index2 == 862 || ((pixel_index2 >= 936) && (pixel_index2 <= 937)) || ((pixel_index2 >= 941) && (pixel_index2 <= 942)) || ((pixel_index2 >= 946) && (pixel_index2 <= 948)) || ((pixel_index2 >= 951) && (pixel_index2 <= 953)) || ((pixel_index2 >= 956) && (pixel_index2 <= 958)) || pixel_index2 == 1034 || pixel_index2 == 1039 || pixel_index2 == 1044 || pixel_index2 == 1046 || pixel_index2 == 1049 || pixel_index2 == 1051 || pixel_index2 == 1054 || ((pixel_index2 >= 1127) && (pixel_index2 <= 1129)) || ((pixel_index2 >= 1132) && (pixel_index2 <= 1134)) || ((pixel_index2 >= 1137) && (pixel_index2 <= 1140)) || ((pixel_index2 >= 1143) && (pixel_index2 <= 1145)) || (pixel_index2 >= 1148) && (pixel_index2 <= 1150)) oled_data2 = 16'b0000011110011110;
            else if (pixel_index2 == 596 || pixel_index2 == 608 || pixel_index2 == 620 || ((pixel_index2 >= 692) && (pixel_index2 <= 693)) || pixel_index2 == 704 || pixel_index2 == 716 || ((pixel_index2 >= 789) && (pixel_index2 <= 790)) || ((pixel_index2 >= 800) && (pixel_index2 <= 801)) || pixel_index2 == 812 || pixel_index2 == 818 || pixel_index2 == 886 || ((pixel_index2 >= 896) && (pixel_index2 <= 897)) || pixel_index2 == 907 || pixel_index2 == 913 || pixel_index2 == 976 || ((pixel_index2 >= 992) && (pixel_index2 <= 993)) || ((pixel_index2 >= 1002) && (pixel_index2 <= 1003)) || pixel_index2 == 1009 || ((pixel_index2 >= 1072) && (pixel_index2 <= 1073)) || pixel_index2 == 1084 || pixel_index2 == 1089 || ((pixel_index2 >= 1097) && (pixel_index2 <= 1099)) || pixel_index2 == 1104 || ((pixel_index2 >= 1168) && (pixel_index2 <= 1170)) || pixel_index2 == 1175 || ((pixel_index2 >= 1180) && (pixel_index2 <= 1181)) || pixel_index2 == 1183 || ((pixel_index2 >= 1185) && (pixel_index2 <= 1186)) || ((pixel_index2 >= 1193) && (pixel_index2 <= 1194)) || ((pixel_index2 >= 1199) && (pixel_index2 <= 1200)) || ((pixel_index2 >= 1265) && (pixel_index2 <= 1267)) || ((pixel_index2 >= 1271) && (pixel_index2 <= 1272)) || ((pixel_index2 >= 1276) && (pixel_index2 <= 1277)) || pixel_index2 == 1279 || ((pixel_index2 >= 1282) && (pixel_index2 <= 1284)) || ((pixel_index2 >= 1288) && (pixel_index2 <= 1290)) || pixel_index2 == 1295 || ((pixel_index2 >= 1362) && (pixel_index2 <= 1365)) || ((pixel_index2 >= 1373) && (pixel_index2 <= 1375)) || ((pixel_index2 >= 1378) && (pixel_index2 <= 1380)) || ((pixel_index2 >= 1384) && (pixel_index2 <= 1386)) || ((pixel_index2 >= 1390) && (pixel_index2 <= 1391)) || ((pixel_index2 >= 1459) && (pixel_index2 <= 1463)) || ((pixel_index2 >= 1470) && (pixel_index2 <= 1471)) || ((pixel_index2 >= 1475) && (pixel_index2 <= 1479)) || pixel_index2 == 1481 || ((pixel_index2 >= 1484) && (pixel_index2 <= 1486)) || pixel_index2 == 1554 || ((pixel_index2 >= 1556) && (pixel_index2 <= 1557)) || pixel_index2 == 1559 || ((pixel_index2 >= 1563) && (pixel_index2 <= 1564)) || pixel_index2 == 1567 || ((pixel_index2 >= 1572) && (pixel_index2 <= 1575)) || pixel_index2 == 1577 || ((pixel_index2 >= 1579) && (pixel_index2 <= 1581)) || pixel_index2 == 1584 || pixel_index2 == 1645 || ((pixel_index2 >= 1650) && (pixel_index2 <= 1651)) || ((pixel_index2 >= 1655) && (pixel_index2 <= 1656)) || ((pixel_index2 >= 1660) && (pixel_index2 <= 1661)) || ((pixel_index2 >= 1676) && (pixel_index2 <= 1677)) || ((pixel_index2 >= 1679) && (pixel_index2 <= 1680)) || pixel_index2 == 1741 || ((pixel_index2 >= 1746) && (pixel_index2 <= 1747)) || ((pixel_index2 >= 1749) && (pixel_index2 <= 1750)) || ((pixel_index2 >= 1752) && (pixel_index2 <= 1753)) || ((pixel_index2 >= 1768) && (pixel_index2 <= 1769)) || pixel_index2 == 1771 || ((pixel_index2 >= 1774) && (pixel_index2 <= 1775)) || ((pixel_index2 >= 1837) && (pixel_index2 <= 1838)) || ((pixel_index2 >= 1843) && (pixel_index2 <= 1846)) || pixel_index2 == 1870 || pixel_index2 == 1934 || ((pixel_index2 >= 1940) && (pixel_index2 <= 1942)) || pixel_index2 == 1965 || pixel_index2 == 1972 || ((pixel_index2 >= 2031) && (pixel_index2 <= 2032)) || ((pixel_index2 >= 2036) && (pixel_index2 <= 2039)) || ((pixel_index2 >= 2059) && (pixel_index2 <= 2060)) || ((pixel_index2 >= 2067) && (pixel_index2 <= 2068)) || ((pixel_index2 >= 2123) && (pixel_index2 <= 2125)) || ((pixel_index2 >= 2128) && (pixel_index2 <= 2130)) || pixel_index2 == 2132 || pixel_index2 == 2135 || ((pixel_index2 >= 2154) && (pixel_index2 <= 2155)) || ((pixel_index2 >= 2162) && (pixel_index2 <= 2164)) || ((pixel_index2 >= 2219) && (pixel_index2 <= 2221)) || ((pixel_index2 >= 2225) && (pixel_index2 <= 2229)) || ((pixel_index2 >= 2249) && (pixel_index2 <= 2250)) || ((pixel_index2 >= 2257) && (pixel_index2 <= 2258)) || ((pixel_index2 >= 2316) && (pixel_index2 <= 2319)) || ((pixel_index2 >= 2323) && (pixel_index2 <= 2326)) || ((pixel_index2 >= 2344) && (pixel_index2 <= 2350)) || ((pixel_index2 >= 2352) && (pixel_index2 <= 2354)) || ((pixel_index2 >= 2415) && (pixel_index2 <= 2416)) || ((pixel_index2 >= 2421) && (pixel_index2 <= 2424)) || ((pixel_index2 >= 2447) && (pixel_index2 <= 2448)) || pixel_index2 == 2520 || ((pixel_index2 >= 2535) && (pixel_index2 <= 2538)) || ((pixel_index2 >= 2541) && (pixel_index2 <= 2543)) || pixel_index2 == 2614 || pixel_index2 == 2627 || ((pixel_index2 >= 2630) && (pixel_index2 <= 2638)) || ((pixel_index2 >= 2707) && (pixel_index2 <= 2712)) || pixel_index2 == 2723 || ((pixel_index2 >= 2726) && (pixel_index2 <= 2727)) || pixel_index2 == 2807 || ((pixel_index2 >= 2810) && (pixel_index2 <= 2811)) || pixel_index2 == 2813 || ((pixel_index2 >= 2819) && (pixel_index2 <= 2822)) || pixel_index2 == 2832 || ((pixel_index2 >= 2902) && (pixel_index2 <= 2903)) || ((pixel_index2 >= 2906) && (pixel_index2 <= 2907)) || pixel_index2 == 2913 || ((pixel_index2 >= 2915) && (pixel_index2 <= 2920)) || pixel_index2 == 2927 || pixel_index2 == 2990 || ((pixel_index2 >= 2997) && (pixel_index2 <= 2998)) || ((pixel_index2 >= 3001) && (pixel_index2 <= 3002)) || ((pixel_index2 >= 3008) && (pixel_index2 <= 3009)) || ((pixel_index2 >= 3022) && (pixel_index2 <= 3023)) || ((pixel_index2 >= 3086) && (pixel_index2 <= 3092)) || ((pixel_index2 >= 3096) && (pixel_index2 <= 3097)) || ((pixel_index2 >= 3105) && (pixel_index2 <= 3107)) || ((pixel_index2 >= 3117) && (pixel_index2 <= 3118)) || ((pixel_index2 >= 3186) && (pixel_index2 <= 3187)) || ((pixel_index2 >= 3203) && (pixel_index2 <= 3213)) || pixel_index2 == 3293 || ((pixel_index2 >= 3301) && (pixel_index2 <= 3306)) || ((pixel_index2 >= 3388) && (pixel_index2 <= 3389)) || pixel_index2 == 3484 || pixel_index2 == 3580) oled_data2 = 16'b0000010100000000;
            else if (pixel_index2 == 1088 || pixel_index2 == 1184 || ((pixel_index2 >= 1280) && (pixel_index2 <= 1281)) || pixel_index2 == 1368 || pixel_index2 == 1372 || ((pixel_index2 >= 1376) && (pixel_index2 <= 1377)) || ((pixel_index2 >= 1464) && (pixel_index2 <= 1465)) || ((pixel_index2 >= 1468) && (pixel_index2 <= 1469)) || ((pixel_index2 >= 1472) && (pixel_index2 <= 1474)) || pixel_index2 == 1480 || pixel_index2 == 1558 || ((pixel_index2 >= 1560) && (pixel_index2 <= 1562)) || ((pixel_index2 >= 1565) && (pixel_index2 <= 1566)) || pixel_index2 == 1568 || pixel_index2 == 1571 || pixel_index2 == 1576 || pixel_index2 == 1654 || ((pixel_index2 >= 1657) && (pixel_index2 <= 1659)) || ((pixel_index2 >= 1662) && (pixel_index2 <= 1664)) || ((pixel_index2 >= 1667) && (pixel_index2 <= 1672)) || ((pixel_index2 >= 1674) && (pixel_index2 <= 1675)) || pixel_index2 == 1751 || ((pixel_index2 >= 1754) && (pixel_index2 <= 1759)) || ((pixel_index2 >= 1763) && (pixel_index2 <= 1767)) || pixel_index2 == 1770 || pixel_index2 == 1773 || ((pixel_index2 >= 1847) && (pixel_index2 <= 1852)) || ((pixel_index2 >= 1860) && (pixel_index2 <= 1869)) || ((pixel_index2 >= 1943) && (pixel_index2 <= 1947)) || ((pixel_index2 >= 1959) && (pixel_index2 <= 1964)) || ((pixel_index2 >= 2040) && (pixel_index2 <= 2041)) || ((pixel_index2 >= 2056) && (pixel_index2 <= 2058)) || ((pixel_index2 >= 2133) && (pixel_index2 <= 2134)) || ((pixel_index2 >= 2136) && (pixel_index2 <= 2137)) || ((pixel_index2 >= 2151) && (pixel_index2 <= 2153)) || ((pixel_index2 >= 2230) && (pixel_index2 <= 2234)) || ((pixel_index2 >= 2245) && (pixel_index2 <= 2248)) || ((pixel_index2 >= 2327) && (pixel_index2 <= 2329)) || pixel_index2 == 2339 || ((pixel_index2 >= 2342) && (pixel_index2 <= 2343)) || ((pixel_index2 >= 2425) && (pixel_index2 <= 2426)) || ((pixel_index2 >= 2434) && (pixel_index2 <= 2446)) || ((pixel_index2 >= 2521) && (pixel_index2 <= 2522)) || ((pixel_index2 >= 2529) && (pixel_index2 <= 2534)) || ((pixel_index2 >= 2539) && (pixel_index2 <= 2540)) || ((pixel_index2 >= 2615) && (pixel_index2 <= 2620)) || ((pixel_index2 >= 2625) && (pixel_index2 <= 2626)) || ((pixel_index2 >= 2628) && (pixel_index2 <= 2629)) || ((pixel_index2 >= 2713) && (pixel_index2 <= 2718)) || ((pixel_index2 >= 2720) && (pixel_index2 <= 2722)) || pixel_index2 == 2725 || pixel_index2 == 2812 || ((pixel_index2 >= 2814) && (pixel_index2 <= 2818)) || ((pixel_index2 >= 2910) && (pixel_index2 <= 2912)) || pixel_index2 == 2914 || ((pixel_index2 >= 3006) && (pixel_index2 <= 3007)) || (pixel_index2 >= 3102) && (pixel_index2 <= 3103)) oled_data2 = 16'b1010011110010100;
            else if (pixel_index2 == 5626 || pixel_index2 == 5630 || ((pixel_index2 >= 5634) && (pixel_index2 <= 5636)) || ((pixel_index2 >= 5638) && (pixel_index2 <= 5641)) || pixel_index2 == 5645 || pixel_index2 == 5649 || pixel_index2 == 5652 || ((pixel_index2 >= 5655) && (pixel_index2 <= 5656)) || ((pixel_index2 >= 5660) && (pixel_index2 <= 5662)) || pixel_index2 == 5729 || pixel_index2 == 5732 || pixel_index2 == 5737 || pixel_index2 == 5741 || pixel_index2 == 5746 || pixel_index2 == 5748 || pixel_index2 == 5750 || pixel_index2 == 5753 || pixel_index2 == 5755 || pixel_index2 == 5818 || pixel_index2 == 5822 || pixel_index2 == 5825 || pixel_index2 == 5828 || ((pixel_index2 >= 5831) && (pixel_index2 <= 5833)) || pixel_index2 == 5837 || ((pixel_index2 >= 5842) && (pixel_index2 <= 5844)) || pixel_index2 == 5846 || pixel_index2 == 5849 || ((pixel_index2 >= 5852) && (pixel_index2 <= 5853)) || pixel_index2 == 5914 || pixel_index2 == 5918 || pixel_index2 == 5921 || pixel_index2 == 5924 || pixel_index2 == 5929 || pixel_index2 == 5933 || pixel_index2 == 5937 || pixel_index2 == 5940 || pixel_index2 == 5942 || pixel_index2 == 5945 || pixel_index2 == 5950 || pixel_index2 == 6010 || pixel_index2 == 6014 || ((pixel_index2 >= 6018) && (pixel_index2 <= 6020)) || ((pixel_index2 >= 6022) && (pixel_index2 <= 6025)) || ((pixel_index2 >= 6027) && (pixel_index2 <= 6031)) || ((pixel_index2 >= 6034) && (pixel_index2 <= 6036)) || ((pixel_index2 >= 6039) && (pixel_index2 <= 6040)) || (pixel_index2 >= 6043) && (pixel_index2 <= 6045)) oled_data2 = 16'b0000000000010100;
            else oled_data2 = 0;
            end
            10: begin
            if (((pixel_index2 >= 138) && (pixel_index2 <= 139)) || ((pixel_index2 >= 217) && (pixel_index2 <= 218)) || ((pixel_index2 >= 225) && (pixel_index2 <= 226)) || ((pixel_index2 >= 234) && (pixel_index2 <= 235)) || ((pixel_index2 >= 313) && (pixel_index2 <= 314)) || ((pixel_index2 >= 321) && (pixel_index2 <= 322)) || ((pixel_index2 >= 494) && (pixel_index2 <= 495)) || ((pixel_index2 >= 527) && (pixel_index2 <= 528)) || ((pixel_index2 >= 590) && (pixel_index2 <= 591)) || ((pixel_index2 >= 623) && (pixel_index2 <= 624)) || ((pixel_index2 >= 1065) && (pixel_index2 <= 1066)) || ((pixel_index2 >= 1161) && (pixel_index2 <= 1162)) || ((pixel_index2 >= 1877) && (pixel_index2 <= 1878)) || ((pixel_index2 >= 1973) && (pixel_index2 <= 1974)) || ((pixel_index2 >= 2025) && (pixel_index2 <= 2026)) || ((pixel_index2 >= 2121) && (pixel_index2 <= 2122)) || ((pixel_index2 >= 2833) && (pixel_index2 <= 2834)) || ((pixel_index2 >= 2929) && (pixel_index2 <= 2930)) || ((pixel_index2 >= 3084) && (pixel_index2 <= 3085)) || ((pixel_index2 >= 3180) && (pixel_index2 <= 3181)) || ((pixel_index2 >= 3593) && (pixel_index2 <= 3594)) || ((pixel_index2 >= 3676) && (pixel_index2 <= 3677)) || ((pixel_index2 >= 3689) && (pixel_index2 <= 3690)) || (pixel_index2 >= 3772) && (pixel_index2 <= 3773)) oled_data2 = 16'b1111011110011110;
            else if (pixel_index2 == 168 || ((pixel_index2 >= 172) && (pixel_index2 <= 175)) || ((pixel_index2 >= 178) && (pixel_index2 <= 180)) || ((pixel_index2 >= 182) && (pixel_index2 <= 185)) || pixel_index2 == 187 || pixel_index2 == 190 || pixel_index2 == 264 || pixel_index2 == 271 || pixel_index2 == 273 || pixel_index2 == 281 || pixel_index2 == 284 || pixel_index2 == 286 || pixel_index2 == 360 || ((pixel_index2 >= 365) && (pixel_index2 <= 367)) || ((pixel_index2 >= 370) && (pixel_index2 <= 371)) || ((pixel_index2 >= 375) && (pixel_index2 <= 377)) || ((pixel_index2 >= 380) && (pixel_index2 <= 382)) || pixel_index2 == 456 || pixel_index2 == 463 || pixel_index2 == 468 || pixel_index2 == 473 || pixel_index2 == 475 || pixel_index2 == 478 || ((pixel_index2 >= 550) && (pixel_index2 <= 554)) || ((pixel_index2 >= 556) && (pixel_index2 <= 559)) || ((pixel_index2 >= 561) && (pixel_index2 <= 563)) || ((pixel_index2 >= 566) && (pixel_index2 <= 569)) || ((pixel_index2 >= 572) && (pixel_index2 <= 574)) || ((pixel_index2 >= 744) && (pixel_index2 <= 746)) || ((pixel_index2 >= 749) && (pixel_index2 <= 751)) || ((pixel_index2 >= 753) && (pixel_index2 <= 756)) || pixel_index2 == 758 || pixel_index2 == 761 || pixel_index2 == 766 || pixel_index2 == 839 || pixel_index2 == 844 || pixel_index2 == 852 || pixel_index2 == 855 || pixel_index2 == 857 || pixel_index2 == 862 || ((pixel_index2 >= 936) && (pixel_index2 <= 937)) || ((pixel_index2 >= 941) && (pixel_index2 <= 942)) || ((pixel_index2 >= 946) && (pixel_index2 <= 948)) || ((pixel_index2 >= 951) && (pixel_index2 <= 953)) || ((pixel_index2 >= 956) && (pixel_index2 <= 958)) || pixel_index2 == 1034 || pixel_index2 == 1039 || pixel_index2 == 1044 || pixel_index2 == 1046 || pixel_index2 == 1049 || pixel_index2 == 1051 || pixel_index2 == 1054 || ((pixel_index2 >= 1127) && (pixel_index2 <= 1129)) || ((pixel_index2 >= 1132) && (pixel_index2 <= 1134)) || ((pixel_index2 >= 1137) && (pixel_index2 <= 1140)) || ((pixel_index2 >= 1143) && (pixel_index2 <= 1145)) || (pixel_index2 >= 1148) && (pixel_index2 <= 1150)) oled_data2 = 16'b1111010100000000;
            else if (pixel_index2 == 592 || pixel_index2 == 596 || pixel_index2 == 608 || pixel_index2 == 620 || ((pixel_index2 >= 687) && (pixel_index2 <= 688)) || ((pixel_index2 >= 692) && (pixel_index2 <= 693)) || pixel_index2 == 704 || pixel_index2 == 716 || ((pixel_index2 >= 784) && (pixel_index2 <= 785)) || ((pixel_index2 >= 789) && (pixel_index2 <= 790)) || ((pixel_index2 >= 800) && (pixel_index2 <= 801)) || pixel_index2 == 812 || pixel_index2 == 818 || ((pixel_index2 >= 880) && (pixel_index2 <= 881)) || pixel_index2 == 886 || ((pixel_index2 >= 896) && (pixel_index2 <= 897)) || pixel_index2 == 907 || pixel_index2 == 913 || pixel_index2 == 977 || pixel_index2 == 992 || pixel_index2 == 1003 || pixel_index2 == 1009 || pixel_index2 == 1084 || ((pixel_index2 >= 1097) && (pixel_index2 <= 1099)) || pixel_index2 == 1104 || pixel_index2 == 1163 || ((pixel_index2 >= 1168) && (pixel_index2 <= 1169)) || pixel_index2 == 1175 || pixel_index2 == 1180 || pixel_index2 == 1186 || ((pixel_index2 >= 1193) && (pixel_index2 <= 1194)) || ((pixel_index2 >= 1199) && (pixel_index2 <= 1200)) || ((pixel_index2 >= 1258) && (pixel_index2 <= 1259)) || ((pixel_index2 >= 1265) && (pixel_index2 <= 1266)) || ((pixel_index2 >= 1271) && (pixel_index2 <= 1272)) || pixel_index2 == 1276 || ((pixel_index2 >= 1282) && (pixel_index2 <= 1284)) || pixel_index2 == 1290 || pixel_index2 == 1295 || ((pixel_index2 >= 1355) && (pixel_index2 <= 1356)) || ((pixel_index2 >= 1362) && (pixel_index2 <= 1363)) || ((pixel_index2 >= 1379) && (pixel_index2 <= 1380)) || pixel_index2 == 1386 || ((pixel_index2 >= 1390) && (pixel_index2 <= 1391)) || ((pixel_index2 >= 1459) && (pixel_index2 <= 1460)) || pixel_index2 == 1477 || pixel_index2 == 1484 || pixel_index2 == 1486 || pixel_index2 == 1554 || ((pixel_index2 >= 1556) && (pixel_index2 <= 1557)) || pixel_index2 == 1573 || ((pixel_index2 >= 1579) && (pixel_index2 <= 1580)) || pixel_index2 == 1584 || pixel_index2 == 1645 || pixel_index2 == 1650 || pixel_index2 == 1656 || pixel_index2 == 1662 || pixel_index2 == 1675 || ((pixel_index2 >= 1679) && (pixel_index2 <= 1680)) || pixel_index2 == 1741 || ((pixel_index2 >= 1746) && (pixel_index2 <= 1747)) || pixel_index2 == 1767 || ((pixel_index2 >= 1837) && (pixel_index2 <= 1838)) || ((pixel_index2 >= 1843) && (pixel_index2 <= 1845)) || pixel_index2 == 1849 || pixel_index2 == 1855 || pixel_index2 == 1870 || pixel_index2 == 1934 || pixel_index2 == 1940 || ((pixel_index2 >= 1950) && (pixel_index2 <= 1951)) || ((pixel_index2 >= 1953) && (pixel_index2 <= 1955)) || pixel_index2 == 1957 || pixel_index2 == 1965 || pixel_index2 == 1972 || ((pixel_index2 >= 2031) && (pixel_index2 <= 2032)) || pixel_index2 == 2036 || pixel_index2 == 2044 || ((pixel_index2 >= 2046) && (pixel_index2 <= 2050)) || ((pixel_index2 >= 2067) && (pixel_index2 <= 2068)) || pixel_index2 == 2123 || ((pixel_index2 >= 2128) && (pixel_index2 <= 2130)) || ((pixel_index2 >= 2139) && (pixel_index2 <= 2145)) || pixel_index2 == 2163 || ((pixel_index2 >= 2218) && (pixel_index2 <= 2220)) || ((pixel_index2 >= 2225) && (pixel_index2 <= 2227)) || ((pixel_index2 >= 2235) && (pixel_index2 <= 2241)) || pixel_index2 == 2250 || ((pixel_index2 >= 2315) && (pixel_index2 <= 2317)) || ((pixel_index2 >= 2323) && (pixel_index2 <= 2324)) || ((pixel_index2 >= 2332) && (pixel_index2 <= 2335)) || pixel_index2 == 2337 || pixel_index2 == 2341 || ((pixel_index2 >= 2345) && (pixel_index2 <= 2346)) || pixel_index2 == 2352 || ((pixel_index2 >= 2413) && (pixel_index2 <= 2414)) || pixel_index2 == 2421 || pixel_index2 == 2424 || ((pixel_index2 >= 2428) && (pixel_index2 <= 2434)) || pixel_index2 == 2447 || pixel_index2 == 2522 || ((pixel_index2 >= 2524) && (pixel_index2 <= 2525)) || ((pixel_index2 >= 2527) && (pixel_index2 <= 2530)) || ((pixel_index2 >= 2542) && (pixel_index2 <= 2543)) || pixel_index2 == 2620 || ((pixel_index2 >= 2623) && (pixel_index2 <= 2624)) || ((pixel_index2 >= 2634) && (pixel_index2 <= 2637)) || pixel_index2 == 2719 || pixel_index2 == 2723 || pixel_index2 == 2727 || ((pixel_index2 >= 2821) && (pixel_index2 <= 2822)) || pixel_index2 == 2832 || ((pixel_index2 >= 2902) && (pixel_index2 <= 2903)) || pixel_index2 == 2910 || ((pixel_index2 >= 2919) && (pixel_index2 <= 2920)) || pixel_index2 == 2927 || pixel_index2 == 2990 || ((pixel_index2 >= 2997) && (pixel_index2 <= 2998)) || ((pixel_index2 >= 3001) && (pixel_index2 <= 3002)) || ((pixel_index2 >= 3022) && (pixel_index2 <= 3023)) || ((pixel_index2 >= 3086) && (pixel_index2 <= 3092)) || ((pixel_index2 >= 3096) && (pixel_index2 <= 3097)) || ((pixel_index2 >= 3102) && (pixel_index2 <= 3103)) || ((pixel_index2 >= 3105) && (pixel_index2 <= 3107)) || ((pixel_index2 >= 3117) && (pixel_index2 <= 3118)) || ((pixel_index2 >= 3186) && (pixel_index2 <= 3187)) || ((pixel_index2 >= 3203) && (pixel_index2 <= 3205)) || pixel_index2 == 3207 || ((pixel_index2 >= 3212) && (pixel_index2 <= 3213)) || pixel_index2 == 3293 || ((pixel_index2 >= 3301) && (pixel_index2 <= 3304)) || ((pixel_index2 >= 3388) && (pixel_index2 <= 3389)) || pixel_index2 == 3484 || pixel_index2 == 3580 || pixel_index2 == 5626 || pixel_index2 == 5630 || ((pixel_index2 >= 5634) && (pixel_index2 <= 5636)) || ((pixel_index2 >= 5638) && (pixel_index2 <= 5641)) || pixel_index2 == 5645 || pixel_index2 == 5649 || pixel_index2 == 5652 || ((pixel_index2 >= 5655) && (pixel_index2 <= 5656)) || ((pixel_index2 >= 5660) && (pixel_index2 <= 5662)) || pixel_index2 == 5729 || pixel_index2 == 5732 || pixel_index2 == 5737 || pixel_index2 == 5741 || pixel_index2 == 5746 || pixel_index2 == 5748 || pixel_index2 == 5750 || pixel_index2 == 5753 || pixel_index2 == 5755 || pixel_index2 == 5818 || pixel_index2 == 5822 || pixel_index2 == 5825 || pixel_index2 == 5828 || ((pixel_index2 >= 5831) && (pixel_index2 <= 5833)) || pixel_index2 == 5837 || ((pixel_index2 >= 5842) && (pixel_index2 <= 5844)) || pixel_index2 == 5846 || pixel_index2 == 5849 || ((pixel_index2 >= 5852) && (pixel_index2 <= 5853)) || pixel_index2 == 5914 || pixel_index2 == 5918 || pixel_index2 == 5921 || pixel_index2 == 5924 || pixel_index2 == 5929 || pixel_index2 == 5933 || pixel_index2 == 5937 || pixel_index2 == 5940 || pixel_index2 == 5942 || pixel_index2 == 5945 || pixel_index2 == 5950 || pixel_index2 == 6010 || pixel_index2 == 6014 || ((pixel_index2 >= 6018) && (pixel_index2 <= 6020)) || ((pixel_index2 >= 6022) && (pixel_index2 <= 6025)) || ((pixel_index2 >= 6027) && (pixel_index2 <= 6031)) || ((pixel_index2 >= 6034) && (pixel_index2 <= 6036)) || ((pixel_index2 >= 6039) && (pixel_index2 <= 6040)) || (pixel_index2 >= 6043) && (pixel_index2 <= 6045)) oled_data2 = 16'b0000010100000000;
            else oled_data2 = 0;
            end
            11: begin
            if (((pixel_index2 >= 49) && (pixel_index2 <= 53)) || (pixel_index2 >= 148) && (pixel_index2 <= 149)) oled_data2 = 16'b1111001010000000;
            else if (((pixel_index2 >= 145) && (pixel_index2 <= 147)) || pixel_index2 == 235 || ((pixel_index2 >= 241) && (pixel_index2 <= 244)) || pixel_index2 == 313 || pixel_index2 == 321 || ((pixel_index2 >= 337) && (pixel_index2 <= 340)) || ((pixel_index2 >= 434) && (pixel_index2 <= 435)) || pixel_index2 == 591 || pixel_index2 == 623 || pixel_index2 == 1162 || pixel_index2 == 1973 || pixel_index2 == 2122 || pixel_index2 == 2833 || pixel_index2 == 3085 || pixel_index2 == 3593 || pixel_index2 == 3676) oled_data2 = 16'b1111011110011110;
            else if (pixel_index2 == 168 || ((pixel_index2 >= 172) && (pixel_index2 <= 175)) || ((pixel_index2 >= 178) && (pixel_index2 <= 180)) || ((pixel_index2 >= 182) && (pixel_index2 <= 185)) || pixel_index2 == 187 || pixel_index2 == 190 || pixel_index2 == 264 || pixel_index2 == 271 || pixel_index2 == 273 || pixel_index2 == 281 || pixel_index2 == 284 || pixel_index2 == 286 || pixel_index2 == 360 || ((pixel_index2 >= 365) && (pixel_index2 <= 367)) || ((pixel_index2 >= 370) && (pixel_index2 <= 371)) || ((pixel_index2 >= 375) && (pixel_index2 <= 377)) || ((pixel_index2 >= 380) && (pixel_index2 <= 382)) || pixel_index2 == 456 || pixel_index2 == 463 || pixel_index2 == 468 || pixel_index2 == 473 || pixel_index2 == 475 || pixel_index2 == 478 || ((pixel_index2 >= 550) && (pixel_index2 <= 554)) || ((pixel_index2 >= 556) && (pixel_index2 <= 559)) || ((pixel_index2 >= 561) && (pixel_index2 <= 563)) || ((pixel_index2 >= 566) && (pixel_index2 <= 569)) || (pixel_index2 >= 572) && (pixel_index2 <= 574)) oled_data2 = 16'b1111000000001010;
            else if (pixel_index2 == 331 || pixel_index2 == 409 || pixel_index2 == 417 || pixel_index2 == 427 || pixel_index2 == 687 || pixel_index2 == 692 || pixel_index2 == 704 || pixel_index2 == 719 || pixel_index2 == 800 || pixel_index2 == 815 || pixel_index2 == 891 || pixel_index2 == 987 || pixel_index2 == 1009 || pixel_index2 == 1098 || pixel_index2 == 1168 || ((pixel_index2 >= 1258) && (pixel_index2 <= 1259)) || pixel_index2 == 1295 || ((pixel_index2 >= 1459) && (pixel_index2 <= 1460)) || pixel_index2 == 1972 || pixel_index2 == 2067 || ((pixel_index2 >= 2218) && (pixel_index2 <= 2219)) || pixel_index2 == 2542 || ((pixel_index2 >= 2637) && (pixel_index2 <= 2638)) || pixel_index2 == 2832 || pixel_index2 == 2901 || ((pixel_index2 >= 2927) && (pixel_index2 <= 2928)) || ((pixel_index2 >= 2990) && (pixel_index2 <= 2991)) || pixel_index2 == 3086 || pixel_index2 == 3091 || pixel_index2 == 3106 || pixel_index2 == 3204 || pixel_index2 == 3304 || pixel_index2 == 3388 || ((pixel_index2 >= 3400) && (pixel_index2 <= 3401)) || pixel_index2 == 3484 || ((pixel_index2 >= 3496) && (pixel_index2 <= 3497)) || (pixel_index2 >= 3580) && (pixel_index2 <= 3581)) oled_data2 = 16'b0000010100000000;
            else if (((pixel_index2 >= 744) && (pixel_index2 <= 746)) || ((pixel_index2 >= 749) && (pixel_index2 <= 751)) || ((pixel_index2 >= 753) && (pixel_index2 <= 756)) || pixel_index2 == 758 || pixel_index2 == 761 || pixel_index2 == 766 || pixel_index2 == 839 || pixel_index2 == 844 || pixel_index2 == 852 || pixel_index2 == 855 || pixel_index2 == 857 || pixel_index2 == 862 || ((pixel_index2 >= 936) && (pixel_index2 <= 937)) || ((pixel_index2 >= 941) && (pixel_index2 <= 942)) || ((pixel_index2 >= 946) && (pixel_index2 <= 948)) || ((pixel_index2 >= 951) && (pixel_index2 <= 953)) || ((pixel_index2 >= 956) && (pixel_index2 <= 958)) || pixel_index2 == 1034 || pixel_index2 == 1039 || pixel_index2 == 1044 || pixel_index2 == 1046 || pixel_index2 == 1049 || pixel_index2 == 1051 || pixel_index2 == 1054 || ((pixel_index2 >= 1127) && (pixel_index2 <= 1129)) || ((pixel_index2 >= 1132) && (pixel_index2 <= 1134)) || ((pixel_index2 >= 1137) && (pixel_index2 <= 1140)) || ((pixel_index2 >= 1143) && (pixel_index2 <= 1145)) || (pixel_index2 >= 1148) && (pixel_index2 <= 1150)) oled_data2 = 16'b1111000000010100;
            else if (pixel_index2 == 5626 || pixel_index2 == 5630 || ((pixel_index2 >= 5634) && (pixel_index2 <= 5636)) || ((pixel_index2 >= 5638) && (pixel_index2 <= 5641)) || pixel_index2 == 5645 || pixel_index2 == 5649 || pixel_index2 == 5652 || ((pixel_index2 >= 5655) && (pixel_index2 <= 5656)) || ((pixel_index2 >= 5660) && (pixel_index2 <= 5662)) || pixel_index2 == 5729 || pixel_index2 == 5732 || pixel_index2 == 5737 || pixel_index2 == 5741 || pixel_index2 == 5746 || pixel_index2 == 5748 || pixel_index2 == 5750 || pixel_index2 == 5753 || pixel_index2 == 5755 || pixel_index2 == 5818 || pixel_index2 == 5822 || pixel_index2 == 5825 || pixel_index2 == 5828 || ((pixel_index2 >= 5831) && (pixel_index2 <= 5833)) || pixel_index2 == 5837 || ((pixel_index2 >= 5842) && (pixel_index2 <= 5844)) || pixel_index2 == 5846 || pixel_index2 == 5849 || ((pixel_index2 >= 5852) && (pixel_index2 <= 5853)) || pixel_index2 == 5914 || pixel_index2 == 5918 || pixel_index2 == 5921 || pixel_index2 == 5924 || pixel_index2 == 5929 || pixel_index2 == 5933 || pixel_index2 == 5937 || pixel_index2 == 5940 || pixel_index2 == 5942 || pixel_index2 == 5945 || pixel_index2 == 5950 || pixel_index2 == 6010 || pixel_index2 == 6014 || ((pixel_index2 >= 6018) && (pixel_index2 <= 6020)) || ((pixel_index2 >= 6022) && (pixel_index2 <= 6025)) || ((pixel_index2 >= 6027) && (pixel_index2 <= 6031)) || ((pixel_index2 >= 6034) && (pixel_index2 <= 6036)) || ((pixel_index2 >= 6039) && (pixel_index2 <= 6040)) || (pixel_index2 >= 6043) && (pixel_index2 <= 6045)) oled_data2 = 16'b1010000000000000;
            else oled_data2 = 0;
            end
            12: begin
            if (pixel_index2 == 168 || ((pixel_index2 >= 172) && (pixel_index2 <= 175)) || ((pixel_index2 >= 178) && (pixel_index2 <= 180)) || ((pixel_index2 >= 182) && (pixel_index2 <= 185)) || pixel_index2 == 187 || pixel_index2 == 190 || pixel_index2 == 264 || pixel_index2 == 271 || pixel_index2 == 273 || pixel_index2 == 281 || pixel_index2 == 284 || pixel_index2 == 286 || pixel_index2 == 360 || ((pixel_index2 >= 365) && (pixel_index2 <= 367)) || ((pixel_index2 >= 370) && (pixel_index2 <= 371)) || ((pixel_index2 >= 375) && (pixel_index2 <= 377)) || ((pixel_index2 >= 380) && (pixel_index2 <= 382)) || pixel_index2 == 456 || pixel_index2 == 463 || pixel_index2 == 468 || pixel_index2 == 473 || pixel_index2 == 475 || pixel_index2 == 478 || ((pixel_index2 >= 550) && (pixel_index2 <= 554)) || ((pixel_index2 >= 556) && (pixel_index2 <= 559)) || ((pixel_index2 >= 561) && (pixel_index2 <= 563)) || ((pixel_index2 >= 566) && (pixel_index2 <= 569)) || ((pixel_index2 >= 572) && (pixel_index2 <= 574)) || ((pixel_index2 >= 744) && (pixel_index2 <= 746)) || ((pixel_index2 >= 749) && (pixel_index2 <= 751)) || ((pixel_index2 >= 753) && (pixel_index2 <= 756)) || pixel_index2 == 758 || pixel_index2 == 761 || pixel_index2 == 766 || pixel_index2 == 839 || pixel_index2 == 844 || pixel_index2 == 852 || pixel_index2 == 855 || pixel_index2 == 857 || pixel_index2 == 862 || ((pixel_index2 >= 936) && (pixel_index2 <= 937)) || ((pixel_index2 >= 941) && (pixel_index2 <= 942)) || ((pixel_index2 >= 946) && (pixel_index2 <= 948)) || ((pixel_index2 >= 951) && (pixel_index2 <= 953)) || ((pixel_index2 >= 956) && (pixel_index2 <= 958)) || pixel_index2 == 1034 || pixel_index2 == 1039 || pixel_index2 == 1044 || pixel_index2 == 1046 || pixel_index2 == 1049 || pixel_index2 == 1051 || pixel_index2 == 1054 || ((pixel_index2 >= 1127) && (pixel_index2 <= 1129)) || ((pixel_index2 >= 1132) && (pixel_index2 <= 1134)) || ((pixel_index2 >= 1137) && (pixel_index2 <= 1140)) || ((pixel_index2 >= 1143) && (pixel_index2 <= 1145)) || (pixel_index2 >= 1148) && (pixel_index2 <= 1150)) oled_data2 = 16'b0000011110011110;
            else if (pixel_index2 == 721 || pixel_index2 == 817 || pixel_index2 == 913 || pixel_index2 == 1009 || pixel_index2 == 1105 || pixel_index2 == 1390 || pixel_index2 == 1486 || pixel_index2 == 1489 || pixel_index2 == 1582 || pixel_index2 == 1585 || pixel_index2 == 1678 || pixel_index2 == 1681 || ((pixel_index2 >= 1773) && (pixel_index2 <= 1775)) || ((pixel_index2 >= 1869) && (pixel_index2 <= 1871)) || pixel_index2 == 1873 || ((pixel_index2 >= 1965) && (pixel_index2 <= 1966)) || ((pixel_index2 >= 2060) && (pixel_index2 <= 2062)) || ((pixel_index2 >= 2156) && (pixel_index2 <= 2158)) || pixel_index2 == 2252 || pixel_index2 == 2254 || ((pixel_index2 >= 2347) && (pixel_index2 <= 2349)) || pixel_index2 == 2443 || pixel_index2 == 2445 || ((pixel_index2 >= 2538) && (pixel_index2 <= 2540)) || ((pixel_index2 >= 2633) && (pixel_index2 <= 2636)) || ((pixel_index2 >= 2729) && (pixel_index2 <= 2731)) || ((pixel_index2 >= 2824) && (pixel_index2 <= 2827)) || ((pixel_index2 >= 2919) && (pixel_index2 <= 2923)) || ((pixel_index2 >= 3014) && (pixel_index2 <= 3015)) || ((pixel_index2 >= 3017) && (pixel_index2 <= 3019)) || ((pixel_index2 >= 3110) && (pixel_index2 <= 3114)) || ((pixel_index2 >= 3207) && (pixel_index2 <= 3210)) || pixel_index2 == 3305 || pixel_index2 == 3401) oled_data2 = 16'b1111001010000000;
            else if (pixel_index2 == 3206 || ((pixel_index2 >= 3301) && (pixel_index2 <= 3303)) || ((pixel_index2 >= 3396) && (pixel_index2 <= 3400)) || ((pixel_index2 >= 3492) && (pixel_index2 <= 3496)) || (pixel_index2 >= 3589) && (pixel_index2 <= 3592)) oled_data2 = 16'b1111011110011110;
            else if (pixel_index2 == 5626 || pixel_index2 == 5630 || ((pixel_index2 >= 5634) && (pixel_index2 <= 5636)) || ((pixel_index2 >= 5638) && (pixel_index2 <= 5641)) || pixel_index2 == 5645 || pixel_index2 == 5649 || pixel_index2 == 5652 || ((pixel_index2 >= 5655) && (pixel_index2 <= 5656)) || ((pixel_index2 >= 5660) && (pixel_index2 <= 5662)) || pixel_index2 == 5729 || pixel_index2 == 5732 || pixel_index2 == 5737 || pixel_index2 == 5741 || pixel_index2 == 5746 || pixel_index2 == 5748 || pixel_index2 == 5750 || pixel_index2 == 5753 || pixel_index2 == 5755 || pixel_index2 == 5818 || pixel_index2 == 5822 || pixel_index2 == 5825 || pixel_index2 == 5828 || ((pixel_index2 >= 5831) && (pixel_index2 <= 5833)) || pixel_index2 == 5837 || ((pixel_index2 >= 5842) && (pixel_index2 <= 5844)) || pixel_index2 == 5846 || pixel_index2 == 5849 || ((pixel_index2 >= 5852) && (pixel_index2 <= 5853)) || pixel_index2 == 5914 || pixel_index2 == 5918 || pixel_index2 == 5921 || pixel_index2 == 5924 || pixel_index2 == 5929 || pixel_index2 == 5933 || pixel_index2 == 5937 || pixel_index2 == 5940 || pixel_index2 == 5942 || pixel_index2 == 5945 || pixel_index2 == 5950 || pixel_index2 == 6010 || pixel_index2 == 6014 || ((pixel_index2 >= 6018) && (pixel_index2 <= 6020)) || ((pixel_index2 >= 6022) && (pixel_index2 <= 6025)) || ((pixel_index2 >= 6027) && (pixel_index2 <= 6031)) || ((pixel_index2 >= 6034) && (pixel_index2 <= 6036)) || ((pixel_index2 >= 6039) && (pixel_index2 <= 6040)) || (pixel_index2 >= 6043) && (pixel_index2 <= 6045)) oled_data2 = 16'b0000000000010100;
            else oled_data2 = 0;
            end                        
        endcase
    end
    if (sw[10] || sw[11] || sw[12] || sw[13] || sw[14]) begin //meme lol, delete if bitstream too slow
        if (((pixel_index2 >= 0) && (pixel_index2 <= 4)) || ((pixel_index2 >= 7) && (pixel_index2 <= 10)) || ((pixel_index2 >= 13) && (pixel_index2 <= 23)) || ((pixel_index2 >= 27) && (pixel_index2 <= 28)) || pixel_index2 == 96 || pixel_index2 == 108 || pixel_index2 == 118 || ((pixel_index2 >= 120) && (pixel_index2 <= 122)) || pixel_index2 == 125 || ((pixel_index2 >= 131) && (pixel_index2 <= 132)) || ((pixel_index2 >= 153) && (pixel_index2 <= 154)) || ((pixel_index2 >= 161) && (pixel_index2 <= 163)) || ((pixel_index2 >= 168) && (pixel_index2 <= 169)) || ((pixel_index2 >= 188) && (pixel_index2 <= 189)) || pixel_index2 == 192 || ((pixel_index2 >= 197) && (pixel_index2 <= 198)) || pixel_index2 == 203 || pixel_index2 == 205 || pixel_index2 == 208 || pixel_index2 == 217 || pixel_index2 == 221 || pixel_index2 == 225 || pixel_index2 == 228 || pixel_index2 == 234 || pixel_index2 == 242 || pixel_index2 == 247 || pixel_index2 == 249 || pixel_index2 == 258 || pixel_index2 == 262 || pixel_index2 == 265 || pixel_index2 == 267 || pixel_index2 == 274 || pixel_index2 == 276 || ((pixel_index2 >= 292) && (pixel_index2 <= 294)) || pixel_index2 == 299 || pixel_index2 == 304 || pixel_index2 == 309 || pixel_index2 == 317 || pixel_index2 == 321 || pixel_index2 == 330 || pixel_index2 == 341 || pixel_index2 == 346 || pixel_index2 == 348 || pixel_index2 == 358 || pixel_index2 == 360 || pixel_index2 == 366 || pixel_index2 == 370 || pixel_index2 == 372 || pixel_index2 == 385 || pixel_index2 == 388 || pixel_index2 == 395 || pixel_index2 == 405 || ((pixel_index2 >= 410) && (pixel_index2 <= 411)) || pixel_index2 == 417 || pixel_index2 == 426 || pixel_index2 == 431 || ((pixel_index2 >= 443) && (pixel_index2 <= 444)) || ((pixel_index2 >= 451) && (pixel_index2 <= 452)) || pixel_index2 == 454 || pixel_index2 == 456 || ((pixel_index2 >= 458) && (pixel_index2 <= 459)) || pixel_index2 == 466 || pixel_index2 == 468 || pixel_index2 == 486 || pixel_index2 == 495 || pixel_index2 == 497 || pixel_index2 == 499 || pixel_index2 == 501 || pixel_index2 == 513 || pixel_index2 == 522 || pixel_index2 == 531 || pixel_index2 == 535 || pixel_index2 == 550 || pixel_index2 == 553 || pixel_index2 == 562 || pixel_index2 == 564 || pixel_index2 == 582 || pixel_index2 == 587 || pixel_index2 == 591 || pixel_index2 == 597 || pixel_index2 == 603 || pixel_index2 == 609 || pixel_index2 == 618 || pixel_index2 == 625 || pixel_index2 == 632 || pixel_index2 == 635 || pixel_index2 == 644 || pixel_index2 == 647 || pixel_index2 == 659 || ((pixel_index2 >= 683) && (pixel_index2 <= 684)) || pixel_index2 == 687 || pixel_index2 == 693 || pixel_index2 == 697 || ((pixel_index2 >= 701) && (pixel_index2 <= 703)) || pixel_index2 == 705 || pixel_index2 == 714 || pixel_index2 == 729 || pixel_index2 == 732 || pixel_index2 == 738 || pixel_index2 == 750 || pixel_index2 == 754 || ((pixel_index2 >= 756) && (pixel_index2 <= 757)) || ((pixel_index2 >= 772) && (pixel_index2 <= 773)) || pixel_index2 == 780 || ((pixel_index2 >= 791) && (pixel_index2 <= 792)) || ((pixel_index2 >= 796) && (pixel_index2 <= 799)) || pixel_index2 == 801 || pixel_index2 == 810 || ((pixel_index2 >= 823) && (pixel_index2 <= 824)) || pixel_index2 == 826 || pixel_index2 == 828 || ((pixel_index2 >= 832) && (pixel_index2 <= 833)) || ((pixel_index2 >= 837) && (pixel_index2 <= 840)) || pixel_index2 == 850 || pixel_index2 == 852 || ((pixel_index2 >= 869) && (pixel_index2 <= 870)) || pixel_index2 == 876 || pixel_index2 == 882 || ((pixel_index2 >= 892) && (pixel_index2 <= 895)) || pixel_index2 == 897 || pixel_index2 == 919 || pixel_index2 == 924 || ((pixel_index2 >= 933) && (pixel_index2 <= 934)) || ((pixel_index2 >= 941) && (pixel_index2 <= 942)) || pixel_index2 == 946 || ((pixel_index2 >= 948) && (pixel_index2 <= 949)) || pixel_index2 == 966 || pixel_index2 == 972 || pixel_index2 == 974 || pixel_index2 == 978 || pixel_index2 == 983 || ((pixel_index2 >= 989) && (pixel_index2 <= 992)) || pixel_index2 == 1004 || pixel_index2 == 1006 || pixel_index2 == 1024 || pixel_index2 == 1035 || pixel_index2 == 1049 || pixel_index2 == 1062 || ((pixel_index2 >= 1066) && (pixel_index2 <= 1067)) || ((pixel_index2 >= 1084) && (pixel_index2 <= 1088)) || ((pixel_index2 >= 1091) && (pixel_index2 <= 1092)) || pixel_index2 == 1158 || ((pixel_index2 >= 1163) && (pixel_index2 <= 1170)) || ((pixel_index2 >= 1173) && (pixel_index2 <= 1193)) || ((pixel_index2 >= 1254) && (pixel_index2 <= 1255)) || ((pixel_index2 >= 1259) && (pixel_index2 <= 1264)) || ((pixel_index2 >= 1270) && (pixel_index2 <= 1272)) || ((pixel_index2 >= 1276) && (pixel_index2 <= 1290)) || ((pixel_index2 >= 1351) && (pixel_index2 <= 1352)) || ((pixel_index2 >= 1355) && (pixel_index2 <= 1360)) || ((pixel_index2 >= 1366) && (pixel_index2 <= 1368)) || ((pixel_index2 >= 1372) && (pixel_index2 <= 1386)) || ((pixel_index2 >= 1447) && (pixel_index2 <= 1455)) || ((pixel_index2 >= 1462) && (pixel_index2 <= 1464)) || ((pixel_index2 >= 1467) && (pixel_index2 <= 1482)) || ((pixel_index2 >= 1543) && (pixel_index2 <= 1551)) || ((pixel_index2 >= 1558) && (pixel_index2 <= 1560)) || pixel_index2 == 1564 || ((pixel_index2 >= 1566) && (pixel_index2 <= 1578)) || ((pixel_index2 >= 1639) && (pixel_index2 <= 1647)) || ((pixel_index2 >= 1654) && (pixel_index2 <= 1656)) || pixel_index2 == 1660 || ((pixel_index2 >= 1662) && (pixel_index2 <= 1676)) || ((pixel_index2 >= 1735) && (pixel_index2 <= 1743)) || ((pixel_index2 >= 1750) && (pixel_index2 <= 1752)) || ((pixel_index2 >= 1757) && (pixel_index2 <= 1760)) || ((pixel_index2 >= 1764) && (pixel_index2 <= 1773)) || ((pixel_index2 >= 1830) && (pixel_index2 <= 1839)) || ((pixel_index2 >= 1846) && (pixel_index2 <= 1848)) || ((pixel_index2 >= 1855) && (pixel_index2 <= 1857)) || ((pixel_index2 >= 1859) && (pixel_index2 <= 1870)) || ((pixel_index2 >= 1926) && (pixel_index2 <= 1935)) || ((pixel_index2 >= 1942) && (pixel_index2 <= 1945)) || ((pixel_index2 >= 1951) && (pixel_index2 <= 1967)) || pixel_index2 == 1987 || ((pixel_index2 >= 2022) && (pixel_index2 <= 2031)) || ((pixel_index2 >= 2038) && (pixel_index2 <= 2041)) || ((pixel_index2 >= 2048) && (pixel_index2 <= 2065)) || pixel_index2 == 2084 || ((pixel_index2 >= 2118) && (pixel_index2 <= 2120)) || ((pixel_index2 >= 2122) && (pixel_index2 <= 2127)) || ((pixel_index2 >= 2134) && (pixel_index2 <= 2137)) || ((pixel_index2 >= 2147) && (pixel_index2 <= 2162)) || pixel_index2 == 2177 || ((pixel_index2 >= 2179) && (pixel_index2 <= 2185)) || ((pixel_index2 >= 2214) && (pixel_index2 <= 2215)) || ((pixel_index2 >= 2218) && (pixel_index2 <= 2223)) || ((pixel_index2 >= 2231) && (pixel_index2 <= 2234)) || ((pixel_index2 >= 2243) && (pixel_index2 <= 2249)) || ((pixel_index2 >= 2251) && (pixel_index2 <= 2259)) || ((pixel_index2 >= 2273) && (pixel_index2 <= 2283)) || ((pixel_index2 >= 2309) && (pixel_index2 <= 2310)) || ((pixel_index2 >= 2314) && (pixel_index2 <= 2319)) || ((pixel_index2 >= 2327) && (pixel_index2 <= 2330)) || ((pixel_index2 >= 2348) && (pixel_index2 <= 2356)) || ((pixel_index2 >= 2369) && (pixel_index2 <= 2380)) || pixel_index2 == 2405 || ((pixel_index2 >= 2409) && (pixel_index2 <= 2415)) || ((pixel_index2 >= 2424) && (pixel_index2 <= 2427)) || ((pixel_index2 >= 2444) && (pixel_index2 <= 2453)) || ((pixel_index2 >= 2465) && (pixel_index2 <= 2477)) || pixel_index2 == 2501 || ((pixel_index2 >= 2505) && (pixel_index2 <= 2510)) || ((pixel_index2 >= 2520) && (pixel_index2 <= 2525)) || ((pixel_index2 >= 2540) && (pixel_index2 <= 2549)) || ((pixel_index2 >= 2561) && (pixel_index2 <= 2574)) || pixel_index2 == 2597 || ((pixel_index2 >= 2601) && (pixel_index2 <= 2606)) || ((pixel_index2 >= 2616) && (pixel_index2 <= 2622)) || ((pixel_index2 >= 2637) && (pixel_index2 <= 2647)) || ((pixel_index2 >= 2658) && (pixel_index2 <= 2671)) || ((pixel_index2 >= 2692) && (pixel_index2 <= 2693)) || ((pixel_index2 >= 2696) && (pixel_index2 <= 2702)) || ((pixel_index2 >= 2712) && (pixel_index2 <= 2724)) || ((pixel_index2 >= 2732) && (pixel_index2 <= 2742)) || ((pixel_index2 >= 2758) && (pixel_index2 <= 2766)) || pixel_index2 == 2788 || ((pixel_index2 >= 2791) && (pixel_index2 <= 2798)) || ((pixel_index2 >= 2809) && (pixel_index2 <= 2812)) || ((pixel_index2 >= 2816) && (pixel_index2 <= 2821)) || ((pixel_index2 >= 2828) && (pixel_index2 <= 2837)) || ((pixel_index2 >= 2858) && (pixel_index2 <= 2862)) || pixel_index2 == 2884 || ((pixel_index2 >= 2887) && (pixel_index2 <= 2894)) || ((pixel_index2 >= 2915) && (pixel_index2 <= 2917)) || ((pixel_index2 >= 2923) && (pixel_index2 <= 2933)) || pixel_index2 == 2980 || ((pixel_index2 >= 2983) && (pixel_index2 <= 2990)) || ((pixel_index2 >= 3012) && (pixel_index2 <= 3016)) || ((pixel_index2 >= 3020) && (pixel_index2 <= 3029)) || pixel_index2 == 3076 || ((pixel_index2 >= 3080) && (pixel_index2 <= 3087)) || ((pixel_index2 >= 3109) && (pixel_index2 <= 3112)) || ((pixel_index2 >= 3115) && (pixel_index2 <= 3126)) || ((pixel_index2 >= 3172) && (pixel_index2 <= 3173)) || ((pixel_index2 >= 3176) && (pixel_index2 <= 3183)) || ((pixel_index2 >= 3205) && (pixel_index2 <= 3208)) || ((pixel_index2 >= 3210) && (pixel_index2 <= 3222)) || ((pixel_index2 >= 3268) && (pixel_index2 <= 3269)) || ((pixel_index2 >= 3272) && (pixel_index2 <= 3279)) || ((pixel_index2 >= 3301) && (pixel_index2 <= 3318)) || pixel_index2 == 3364 || pixel_index2 == 3369 || ((pixel_index2 >= 3372) && (pixel_index2 <= 3375)) || ((pixel_index2 >= 3398) && (pixel_index2 <= 3415)) || pixel_index2 == 3460 || ((pixel_index2 >= 3469) && (pixel_index2 <= 3471)) || ((pixel_index2 >= 3495) && (pixel_index2 <= 3511)) || pixel_index2 == 3556 || ((pixel_index2 >= 3565) && (pixel_index2 <= 3568)) || ((pixel_index2 >= 3592) && (pixel_index2 <= 3607)) || pixel_index2 == 3652 || ((pixel_index2 >= 3662) && (pixel_index2 <= 3664)) || ((pixel_index2 >= 3690) && (pixel_index2 <= 3704)) || ((pixel_index2 >= 3748) && (pixel_index2 <= 3749)) || ((pixel_index2 >= 3759) && (pixel_index2 <= 3762)) || ((pixel_index2 >= 3788) && (pixel_index2 <= 3801)) || ((pixel_index2 >= 3844) && (pixel_index2 <= 3845)) || ((pixel_index2 >= 3855) && (pixel_index2 <= 3861)) || ((pixel_index2 >= 3885) && (pixel_index2 <= 3897)) || ((pixel_index2 >= 3941) && (pixel_index2 <= 3942)) || ((pixel_index2 >= 3953) && (pixel_index2 <= 3963)) || ((pixel_index2 >= 3982) && (pixel_index2 <= 3995)) || ((pixel_index2 >= 4037) && (pixel_index2 <= 4039)) || ((pixel_index2 >= 4050) && (pixel_index2 <= 4059)) || ((pixel_index2 >= 4079) && (pixel_index2 <= 4094)) || ((pixel_index2 >= 4134) && (pixel_index2 <= 4135)) || ((pixel_index2 >= 4146) && (pixel_index2 <= 4156)) || ((pixel_index2 >= 4176) && (pixel_index2 <= 4191)) || ((pixel_index2 >= 4231) && (pixel_index2 <= 4234)) || ((pixel_index2 >= 4243) && (pixel_index2 <= 4252)) || ((pixel_index2 >= 4259) && (pixel_index2 <= 4260)) || ((pixel_index2 >= 4273) && (pixel_index2 <= 4288)) || pixel_index2 == 4330 || ((pixel_index2 >= 4341) && (pixel_index2 <= 4358)) || ((pixel_index2 >= 4370) && (pixel_index2 <= 4383)) || ((pixel_index2 >= 4426) && (pixel_index2 <= 4428)) || ((pixel_index2 >= 4436) && (pixel_index2 <= 4438)) || ((pixel_index2 >= 4440) && (pixel_index2 <= 4455)) || ((pixel_index2 >= 4466) && (pixel_index2 <= 4477)) || ((pixel_index2 >= 4523) && (pixel_index2 <= 4525)) || ((pixel_index2 >= 4532) && (pixel_index2 <= 4550)) || pixel_index2 == 4552 || ((pixel_index2 >= 4562) && (pixel_index2 <= 4567)) || ((pixel_index2 >= 4621) && (pixel_index2 <= 4646)) || ((pixel_index2 >= 4659) && (pixel_index2 <= 4663)) || ((pixel_index2 >= 4719) && (pixel_index2 <= 4744)) || ((pixel_index2 >= 4750) && (pixel_index2 <= 4752)) || ((pixel_index2 >= 4755) && (pixel_index2 <= 4759)) || ((pixel_index2 >= 4818) && (pixel_index2 <= 4850)) || ((pixel_index2 >= 4852) && (pixel_index2 <= 4854)) || ((pixel_index2 >= 4869) && (pixel_index2 <= 4871)) || ((pixel_index2 >= 4916) && (pixel_index2 <= 4919)) || pixel_index2 == 4924 || pixel_index2 == 4928 || pixel_index2 == 4932 || pixel_index2 == 4938 || ((pixel_index2 >= 4946) && (pixel_index2 <= 4948)) || ((pixel_index2 >= 5013) && (pixel_index2 <= 5015)) || ((pixel_index2 >= 5020) && (pixel_index2 <= 5021)) || pixel_index2 == 5025 || pixel_index2 == 5033 || ((pixel_index2 >= 5042) && (pixel_index2 <= 5043)) || pixel_index2 == 5045 || pixel_index2 == 5057 || ((pixel_index2 >= 5109) && (pixel_index2 <= 5111)) || ((pixel_index2 >= 5116) && (pixel_index2 <= 5117)) || pixel_index2 == 5121 || pixel_index2 == 5124 || pixel_index2 == 5131 || ((pixel_index2 >= 5138) && (pixel_index2 <= 5139)) || pixel_index2 == 5153 || ((pixel_index2 >= 5205) && (pixel_index2 <= 5207)) || ((pixel_index2 >= 5212) && (pixel_index2 <= 5213)) || pixel_index2 == 5217 || pixel_index2 == 5220 || pixel_index2 == 5227 || pixel_index2 == 5229 || ((pixel_index2 >= 5234) && (pixel_index2 <= 5235)) || pixel_index2 == 5242 || pixel_index2 == 5249 || pixel_index2 == 5257 || ((pixel_index2 >= 5300) && (pixel_index2 <= 5303)) || ((pixel_index2 >= 5308) && (pixel_index2 <= 5309)) || pixel_index2 == 5313 || pixel_index2 == 5316 || pixel_index2 == 5323 || pixel_index2 == 5325 || ((pixel_index2 >= 5330) && (pixel_index2 <= 5331)) || pixel_index2 == 5338 || pixel_index2 == 5345 || ((pixel_index2 >= 5353) && (pixel_index2 <= 5354)) || ((pixel_index2 >= 5396) && (pixel_index2 <= 5399)) || ((pixel_index2 >= 5404) && (pixel_index2 <= 5405)) || pixel_index2 == 5412 || pixel_index2 == 5419 || pixel_index2 == 5421 || ((pixel_index2 >= 5426) && (pixel_index2 <= 5427)) || pixel_index2 == 5434 || pixel_index2 == 5436 || pixel_index2 == 5438 || pixel_index2 == 5441 || pixel_index2 == 5445 || ((pixel_index2 >= 5449) && (pixel_index2 <= 5455)) || ((pixel_index2 >= 5493) && (pixel_index2 <= 5495)) || ((pixel_index2 >= 5500) && (pixel_index2 <= 5501)) || pixel_index2 == 5503 || pixel_index2 == 5508 || pixel_index2 == 5515 || pixel_index2 == 5517 || pixel_index2 == 5522 || pixel_index2 == 5530 || pixel_index2 == 5532 || pixel_index2 == 5537 || pixel_index2 == 5539 || ((pixel_index2 >= 5545) && (pixel_index2 <= 5552)) || pixel_index2 == 5597 || ((pixel_index2 >= 5599) && (pixel_index2 <= 5600)) || pixel_index2 == 5604 || pixel_index2 == 5611 || pixel_index2 == 5613 || ((pixel_index2 >= 5618) && (pixel_index2 <= 5619)) || pixel_index2 == 5626 || pixel_index2 == 5633 || ((pixel_index2 >= 5641) && (pixel_index2 <= 5645)) || pixel_index2 == 5693 || ((pixel_index2 >= 5695) && (pixel_index2 <= 5696)) || pixel_index2 == 5700 || pixel_index2 == 5707 || pixel_index2 == 5709 || ((pixel_index2 >= 5714) && (pixel_index2 <= 5715)) || pixel_index2 == 5729 || ((pixel_index2 >= 5788) && (pixel_index2 <= 5789)) || pixel_index2 == 5791 || pixel_index2 == 5799 || pixel_index2 == 5806 || pixel_index2 == 5815 || pixel_index2 == 5822 || pixel_index2 == 5825 || pixel_index2 == 5829 || ((pixel_index2 >= 5879) && (pixel_index2 <= 5887)) || ((pixel_index2 >= 5889) && (pixel_index2 <= 5890)) || pixel_index2 == 5894 || pixel_index2 == 5896 || ((pixel_index2 >= 5901) && (pixel_index2 <= 5904)) || pixel_index2 == 5910 || ((pixel_index2 >= 5917) && (pixel_index2 <= 5920)) || (pixel_index2 >= 5924) && (pixel_index2 <= 5927)) oled_data2 = 16'b1010010100010100;
        else if (((pixel_index2 >= 5) && (pixel_index2 <= 6)) || ((pixel_index2 >= 11) && (pixel_index2 <= 12)) || ((pixel_index2 >= 101) && (pixel_index2 <= 102)) || pixel_index2 == 107 || pixel_index2 == 237 || pixel_index2 == 289 || pixel_index2 == 491 || ((pixel_index2 >= 1159) && (pixel_index2 <= 1162)) || ((pixel_index2 >= 1256) && (pixel_index2 <= 1258)) || ((pixel_index2 >= 1273) && (pixel_index2 <= 1275)) || ((pixel_index2 >= 1353) && (pixel_index2 <= 1354)) || ((pixel_index2 >= 1369) && (pixel_index2 <= 1371)) || ((pixel_index2 >= 1465) && (pixel_index2 <= 1466)) || ((pixel_index2 >= 1561) && (pixel_index2 <= 1563)) || pixel_index2 == 1565 || ((pixel_index2 >= 1657) && (pixel_index2 <= 1659)) || pixel_index2 == 1661 || ((pixel_index2 >= 1753) && (pixel_index2 <= 1756)) || ((pixel_index2 >= 1761) && (pixel_index2 <= 1763)) || ((pixel_index2 >= 1849) && (pixel_index2 <= 1854)) || pixel_index2 == 1858 || ((pixel_index2 >= 1946) && (pixel_index2 <= 1950)) || ((pixel_index2 >= 2042) && (pixel_index2 <= 2047)) || pixel_index2 == 2121 || ((pixel_index2 >= 2138) && (pixel_index2 <= 2146)) || ((pixel_index2 >= 2216) && (pixel_index2 <= 2217)) || ((pixel_index2 >= 2235) && (pixel_index2 <= 2242)) || pixel_index2 == 2250 || ((pixel_index2 >= 2311) && (pixel_index2 <= 2313)) || ((pixel_index2 >= 2331) && (pixel_index2 <= 2347)) || ((pixel_index2 >= 2406) && (pixel_index2 <= 2408)) || ((pixel_index2 >= 2428) && (pixel_index2 <= 2443)) || ((pixel_index2 >= 2502) && (pixel_index2 <= 2504)) || ((pixel_index2 >= 2526) && (pixel_index2 <= 2539)) || ((pixel_index2 >= 2598) && (pixel_index2 <= 2600)) || ((pixel_index2 >= 2623) && (pixel_index2 <= 2636)) || ((pixel_index2 >= 2694) && (pixel_index2 <= 2695)) || ((pixel_index2 >= 2725) && (pixel_index2 <= 2731)) || ((pixel_index2 >= 2789) && (pixel_index2 <= 2790)) || ((pixel_index2 >= 2822) && (pixel_index2 <= 2827)) || ((pixel_index2 >= 2885) && (pixel_index2 <= 2886)) || ((pixel_index2 >= 2918) && (pixel_index2 <= 2922)) || ((pixel_index2 >= 2981) && (pixel_index2 <= 2982)) || ((pixel_index2 >= 3017) && (pixel_index2 <= 3019)) || ((pixel_index2 >= 3077) && (pixel_index2 <= 3079)) || ((pixel_index2 >= 3113) && (pixel_index2 <= 3114)) || ((pixel_index2 >= 3174) && (pixel_index2 <= 3175)) || pixel_index2 == 3209 || ((pixel_index2 >= 3270) && (pixel_index2 <= 3271)) || ((pixel_index2 >= 3365) && (pixel_index2 <= 3368)) || ((pixel_index2 >= 3370) && (pixel_index2 <= 3371)) || ((pixel_index2 >= 3461) && (pixel_index2 <= 3468)) || ((pixel_index2 >= 3557) && (pixel_index2 <= 3564)) || ((pixel_index2 >= 3653) && (pixel_index2 <= 3661)) || ((pixel_index2 >= 3750) && (pixel_index2 <= 3758)) || ((pixel_index2 >= 3846) && (pixel_index2 <= 3854)) || ((pixel_index2 >= 3943) && (pixel_index2 <= 3952)) || ((pixel_index2 >= 4040) && (pixel_index2 <= 4049)) || ((pixel_index2 >= 4136) && (pixel_index2 <= 4145)) || ((pixel_index2 >= 4235) && (pixel_index2 <= 4242)) || ((pixel_index2 >= 4331) && (pixel_index2 <= 4340)) || ((pixel_index2 >= 4429) && (pixel_index2 <= 4435)) || pixel_index2 == 4439 || ((pixel_index2 >= 4526) && (pixel_index2 <= 4531)) || pixel_index2 == 5523) oled_data2 = 16'b1111010100010100;
        else if (pixel_index2 == 24 || ((pixel_index2 >= 32) && (pixel_index2 <= 33)) || ((pixel_index2 >= 38) && (pixel_index2 <= 39)) || pixel_index2 == 98 || ((pixel_index2 >= 109) && (pixel_index2 <= 111)) || ((pixel_index2 >= 115) && (pixel_index2 <= 116)) || ((pixel_index2 >= 127) && (pixel_index2 <= 128)) || ((pixel_index2 >= 136) && (pixel_index2 <= 137)) || pixel_index2 == 142 || pixel_index2 == 144 || pixel_index2 == 176 || pixel_index2 == 224 || pixel_index2 == 695 || pixel_index2 == 1063 || ((pixel_index2 >= 1098) && (pixel_index2 <= 1099)) || pixel_index2 == 1157 || ((pixel_index2 >= 1195) && (pixel_index2 <= 1198)) || pixel_index2 == 1253 || ((pixel_index2 >= 1291) && (pixel_index2 <= 1295)) || ((pixel_index2 >= 1307) && (pixel_index2 <= 1310)) || pixel_index2 == 1334 || ((pixel_index2 >= 1388) && (pixel_index2 <= 1393)) || ((pixel_index2 >= 1404) && (pixel_index2 <= 1407)) || pixel_index2 == 1430 || ((pixel_index2 >= 1484) && (pixel_index2 <= 1492)) || ((pixel_index2 >= 1502) && (pixel_index2 <= 1504)) || ((pixel_index2 >= 1506) && (pixel_index2 <= 1512)) || ((pixel_index2 >= 1582) && (pixel_index2 <= 1591)) || ((pixel_index2 >= 1599) && (pixel_index2 <= 1609)) || ((pixel_index2 >= 1678) && (pixel_index2 <= 1688)) || ((pixel_index2 >= 1695) && (pixel_index2 <= 1705)) || ((pixel_index2 >= 1776) && (pixel_index2 <= 1784)) || ((pixel_index2 >= 1792) && (pixel_index2 <= 1803)) || pixel_index2 == 1816 || ((pixel_index2 >= 1873) && (pixel_index2 <= 1880)) || ((pixel_index2 >= 1887) && (pixel_index2 <= 1889)) || ((pixel_index2 >= 1897) && (pixel_index2 <= 1899)) || ((pixel_index2 >= 1970) && (pixel_index2 <= 1976)) || ((pixel_index2 >= 1983) && (pixel_index2 <= 1984)) || ((pixel_index2 >= 1994) && (pixel_index2 <= 1995)) || ((pixel_index2 >= 2009) && (pixel_index2 <= 2010)) || pixel_index2 == 2021 || ((pixel_index2 >= 2068) && (pixel_index2 <= 2072)) || ((pixel_index2 >= 2079) && (pixel_index2 <= 2080)) || pixel_index2 == 2092 || ((pixel_index2 >= 2104) && (pixel_index2 <= 2106)) || ((pixel_index2 >= 2165) && (pixel_index2 <= 2168)) || ((pixel_index2 >= 2174) && (pixel_index2 <= 2176)) || ((pixel_index2 >= 2189) && (pixel_index2 <= 2190)) || ((pixel_index2 >= 2199) && (pixel_index2 <= 2203)) || ((pixel_index2 >= 2261) && (pixel_index2 <= 2265)) || ((pixel_index2 >= 2270) && (pixel_index2 <= 2271)) || ((pixel_index2 >= 2287) && (pixel_index2 <= 2289)) || ((pixel_index2 >= 2295) && (pixel_index2 <= 2299)) || pixel_index2 == 2308 || ((pixel_index2 >= 2357) && (pixel_index2 <= 2367)) || ((pixel_index2 >= 2384) && (pixel_index2 <= 2386)) || ((pixel_index2 >= 2390) && (pixel_index2 <= 2396)) || pixel_index2 == 2404 || ((pixel_index2 >= 2455) && (pixel_index2 <= 2463)) || ((pixel_index2 >= 2481) && (pixel_index2 <= 2483)) || ((pixel_index2 >= 2486) && (pixel_index2 <= 2492)) || ((pixel_index2 >= 2552) && (pixel_index2 <= 2559)) || ((pixel_index2 >= 2578) && (pixel_index2 <= 2588)) || ((pixel_index2 >= 2649) && (pixel_index2 <= 2654)) || ((pixel_index2 >= 2674) && (pixel_index2 <= 2684)) || ((pixel_index2 >= 2745) && (pixel_index2 <= 2750)) || ((pixel_index2 >= 2770) && (pixel_index2 <= 2780)) || pixel_index2 == 2803 || ((pixel_index2 >= 2848) && (pixel_index2 <= 2854)) || ((pixel_index2 >= 2865) && (pixel_index2 <= 2866)) || ((pixel_index2 >= 2868) && (pixel_index2 <= 2877)) || pixel_index2 == 2883 || ((pixel_index2 >= 2898) && (pixel_index2 <= 2900)) || ((pixel_index2 >= 2911) && (pixel_index2 <= 2913)) || ((pixel_index2 >= 2942) && (pixel_index2 <= 2943)) || ((pixel_index2 >= 2949) && (pixel_index2 <= 2955)) || ((pixel_index2 >= 2960) && (pixel_index2 <= 2962)) || ((pixel_index2 >= 2964) && (pixel_index2 <= 2973)) || pixel_index2 == 2979 || pixel_index2 == 2994 || ((pixel_index2 >= 3009) && (pixel_index2 <= 3010)) || ((pixel_index2 >= 3038) && (pixel_index2 <= 3039)) || ((pixel_index2 >= 3059) && (pixel_index2 <= 3069)) || ((pixel_index2 >= 3106) && (pixel_index2 <= 3107)) || ((pixel_index2 >= 3134) && (pixel_index2 <= 3136)) || ((pixel_index2 >= 3155) && (pixel_index2 <= 3165)) || pixel_index2 == 3171 || pixel_index2 == 3185 || ((pixel_index2 >= 3202) && (pixel_index2 <= 3204)) || ((pixel_index2 >= 3230) && (pixel_index2 <= 3231)) || ((pixel_index2 >= 3251) && (pixel_index2 <= 3261)) || pixel_index2 == 3267 || pixel_index2 == 3281 || ((pixel_index2 >= 3299) && (pixel_index2 <= 3300)) || ((pixel_index2 >= 3326) && (pixel_index2 <= 3327)) || pixel_index2 == 3348 || ((pixel_index2 >= 3351) && (pixel_index2 <= 3357)) || pixel_index2 == 3363 || pixel_index2 == 3377 || ((pixel_index2 >= 3395) && (pixel_index2 <= 3396)) || ((pixel_index2 >= 3422) && (pixel_index2 <= 3423)) || ((pixel_index2 >= 3444) && (pixel_index2 <= 3445)) || ((pixel_index2 >= 3448) && (pixel_index2 <= 3453)) || pixel_index2 == 3459 || pixel_index2 == 3473 || ((pixel_index2 >= 3491) && (pixel_index2 <= 3492)) || ((pixel_index2 >= 3519) && (pixel_index2 <= 3520)) || ((pixel_index2 >= 3541) && (pixel_index2 <= 3542)) || ((pixel_index2 >= 3545) && (pixel_index2 <= 3549)) || pixel_index2 == 3555 || pixel_index2 == 3569 || ((pixel_index2 >= 3586) && (pixel_index2 <= 3589)) || ((pixel_index2 >= 3614) && (pixel_index2 <= 3617)) || ((pixel_index2 >= 3638) && (pixel_index2 <= 3645)) || pixel_index2 == 3651 || ((pixel_index2 >= 3681) && (pixel_index2 <= 3684)) || ((pixel_index2 >= 3710) && (pixel_index2 <= 3714)) || ((pixel_index2 >= 3734) && (pixel_index2 <= 3735)) || pixel_index2 == 3741 || ((pixel_index2 >= 3763) && (pixel_index2 <= 3764)) || ((pixel_index2 >= 3774) && (pixel_index2 <= 3776)) || ((pixel_index2 >= 3778) && (pixel_index2 <= 3779)) || ((pixel_index2 >= 3807) && (pixel_index2 <= 3811)) || pixel_index2 == 3830 || pixel_index2 == 3837 || pixel_index2 == 3872 || ((pixel_index2 >= 3905) && (pixel_index2 <= 3909)) || pixel_index2 == 3926 || pixel_index2 == 3933 || pixel_index2 == 3939 || ((pixel_index2 >= 4002) && (pixel_index2 <= 4007)) || ((pixel_index2 >= 4019) && (pixel_index2 <= 4021)) || pixel_index2 == 4035 || ((pixel_index2 >= 4100) && (pixel_index2 <= 4117)) || pixel_index2 == 4131 || ((pixel_index2 >= 4196) && (pixel_index2 <= 4213)) || pixel_index2 == 4220 || ((pixel_index2 >= 4227) && (pixel_index2 <= 4228)) || ((pixel_index2 >= 4293) && (pixel_index2 <= 4300)) || ((pixel_index2 >= 4302) && (pixel_index2 <= 4309)) || ((pixel_index2 >= 4323) && (pixel_index2 <= 4324)) || ((pixel_index2 >= 4398) && (pixel_index2 <= 4404)) || pixel_index2 == 4419 || ((pixel_index2 >= 4495) && (pixel_index2 <= 4499)) || pixel_index2 == 4504 || ((pixel_index2 >= 4506) && (pixel_index2 <= 4508)) || ((pixel_index2 >= 4514) && (pixel_index2 <= 4515)) || pixel_index2 == 4520 || ((pixel_index2 >= 4592) && (pixel_index2 <= 4595)) || ((pixel_index2 >= 4599) && (pixel_index2 <= 4605)) || pixel_index2 == 4610 || ((pixel_index2 >= 4616) && (pixel_index2 <= 4617)) || ((pixel_index2 >= 4688) && (pixel_index2 <= 4692)) || ((pixel_index2 >= 4695) && (pixel_index2 <= 4698)) || ((pixel_index2 >= 4700) && (pixel_index2 <= 4701)) || pixel_index2 == 4706 || ((pixel_index2 >= 4712) && (pixel_index2 <= 4715)) || ((pixel_index2 >= 4785) && (pixel_index2 <= 4792)) || ((pixel_index2 >= 4796) && (pixel_index2 <= 4797)) || pixel_index2 == 4802 || ((pixel_index2 >= 4809) && (pixel_index2 <= 4811)) || ((pixel_index2 >= 4880) && (pixel_index2 <= 4884)) || ((pixel_index2 >= 4892) && (pixel_index2 <= 4893)) || pixel_index2 == 4898 || ((pixel_index2 >= 4907) && (pixel_index2 <= 4910)) || pixel_index2 == 4931 || pixel_index2 == 4937 || ((pixel_index2 >= 4975) && (pixel_index2 <= 4977)) || ((pixel_index2 >= 4987) && (pixel_index2 <= 4989)) || ((pixel_index2 >= 4994) && (pixel_index2 <= 4995)) || ((pixel_index2 >= 5001) && (pixel_index2 <= 5009)) || ((pixel_index2 >= 5070) && (pixel_index2 <= 5073)) || ((pixel_index2 >= 5082) && (pixel_index2 <= 5085)) || ((pixel_index2 >= 5090) && (pixel_index2 <= 5091)) || ((pixel_index2 >= 5097) && (pixel_index2 <= 5105)) || ((pixel_index2 >= 5166) && (pixel_index2 <= 5169)) || ((pixel_index2 >= 5175) && (pixel_index2 <= 5182)) || pixel_index2 == 5187 || ((pixel_index2 >= 5193) && (pixel_index2 <= 5201)) || ((pixel_index2 >= 5261) && (pixel_index2 <= 5266)) || ((pixel_index2 >= 5271) && (pixel_index2 <= 5278)) || pixel_index2 == 5283 || ((pixel_index2 >= 5289) && (pixel_index2 <= 5296)) || pixel_index2 == 5361 || ((pixel_index2 >= 5363) && (pixel_index2 <= 5374)) || pixel_index2 == 5378 || ((pixel_index2 >= 5384) && (pixel_index2 <= 5392)) || ((pixel_index2 >= 5465) && (pixel_index2 <= 5470)) || pixel_index2 == 5474 || ((pixel_index2 >= 5479) && (pixel_index2 <= 5490)) || ((pixel_index2 >= 5561) && (pixel_index2 <= 5568)) || ((pixel_index2 >= 5573) && (pixel_index2 <= 5581)) || pixel_index2 == 5661 || pixel_index2 == 5663 || ((pixel_index2 >= 5669) && (pixel_index2 <= 5673)) || pixel_index2 == 5736 || ((pixel_index2 >= 5739) && (pixel_index2 <= 5740)) || pixel_index2 == 5747 || pixel_index2 == 5759 || ((pixel_index2 >= 5764) && (pixel_index2 <= 5767)) || ((pixel_index2 >= 5844) && (pixel_index2 <= 5845)) || pixel_index2 == 5855 || ((pixel_index2 >= 5859) && (pixel_index2 <= 5861)) || ((pixel_index2 >= 5945) && (pixel_index2 <= 5946)) || pixel_index2 == 5951 || ((pixel_index2 >= 5954) && (pixel_index2 <= 5955)) || pixel_index2 == 6044 || pixel_index2 == 6047 || pixel_index2 == 6050 || (pixel_index2 >= 6142) && (pixel_index2 <= 6143)) oled_data2 = 16'b1010001010001010;
        else if (((pixel_index2 >= 25) && (pixel_index2 <= 26)) || ((pixel_index2 >= 34) && (pixel_index2 <= 37)) || ((pixel_index2 >= 40) && (pixel_index2 <= 95)) || pixel_index2 == 97 || pixel_index2 == 100 || pixel_index2 == 103 || pixel_index2 == 106 || ((pixel_index2 >= 112) && (pixel_index2 <= 113)) || pixel_index2 == 117 || pixel_index2 == 119 || pixel_index2 == 123 || ((pixel_index2 >= 129) && (pixel_index2 <= 130)) || ((pixel_index2 >= 133) && (pixel_index2 <= 135)) || ((pixel_index2 >= 138) && (pixel_index2 <= 141)) || pixel_index2 == 143 || ((pixel_index2 >= 145) && (pixel_index2 <= 148)) || ((pixel_index2 >= 150) && (pixel_index2 <= 151)) || pixel_index2 == 155 || ((pixel_index2 >= 157) && (pixel_index2 <= 160)) || ((pixel_index2 >= 164) && (pixel_index2 <= 167)) || ((pixel_index2 >= 171) && (pixel_index2 <= 175)) || ((pixel_index2 >= 178) && (pixel_index2 <= 187)) || ((pixel_index2 >= 190) && (pixel_index2 <= 191)) || pixel_index2 == 193 || pixel_index2 == 196 || pixel_index2 == 199 || pixel_index2 == 209 || ((pixel_index2 >= 213) && (pixel_index2 <= 214)) || ((pixel_index2 >= 235) && (pixel_index2 <= 236)) || pixel_index2 == 245 || ((pixel_index2 >= 252) && (pixel_index2 <= 255)) || pixel_index2 == 268 || pixel_index2 == 277 || ((pixel_index2 >= 281) && (pixel_index2 <= 282)) || pixel_index2 == 286 || pixel_index2 == 288 || pixel_index2 == 300 || pixel_index2 == 305 || pixel_index2 == 310 || pixel_index2 == 316 || pixel_index2 == 320 || ((pixel_index2 >= 323) && (pixel_index2 <= 324)) || ((pixel_index2 >= 331) && (pixel_index2 <= 332)) || pixel_index2 == 345 || ((pixel_index2 >= 349) && (pixel_index2 <= 351)) || pixel_index2 == 357 || pixel_index2 == 361 || ((pixel_index2 >= 364) && (pixel_index2 <= 365)) || pixel_index2 == 373 || ((pixel_index2 >= 377) && (pixel_index2 <= 378)) || pixel_index2 == 382 || pixel_index2 == 384 || pixel_index2 == 396 || pixel_index2 == 401 || pixel_index2 == 406 || ((pixel_index2 >= 412) && (pixel_index2 <= 415)) || pixel_index2 == 419 || ((pixel_index2 >= 427) && (pixel_index2 <= 428)) || ((pixel_index2 >= 441) && (pixel_index2 <= 442)) || ((pixel_index2 >= 445) && (pixel_index2 <= 447)) || pixel_index2 == 457 || ((pixel_index2 >= 460) && (pixel_index2 <= 462)) || pixel_index2 == 469 || ((pixel_index2 >= 473) && (pixel_index2 <= 474)) || pixel_index2 == 478 || pixel_index2 == 481 || pixel_index2 == 490 || pixel_index2 == 492 || pixel_index2 == 502 || ((pixel_index2 >= 506) && (pixel_index2 <= 508)) || pixel_index2 == 515 || ((pixel_index2 >= 523) && (pixel_index2 <= 524)) || pixel_index2 == 527 || pixel_index2 == 538 || ((pixel_index2 >= 541) && (pixel_index2 <= 543)) || pixel_index2 == 547 || pixel_index2 == 549 || ((pixel_index2 >= 555) && (pixel_index2 <= 558)) || pixel_index2 == 565 || ((pixel_index2 >= 570) && (pixel_index2 <= 571)) || pixel_index2 == 574 || ((pixel_index2 >= 576) && (pixel_index2 <= 577)) || pixel_index2 == 580 || pixel_index2 == 583 || pixel_index2 == 586 || pixel_index2 == 588 || pixel_index2 == 595 || ((pixel_index2 >= 598) && (pixel_index2 <= 599)) || ((pixel_index2 >= 604) && (pixel_index2 <= 607)) || pixel_index2 == 611 || ((pixel_index2 >= 619) && (pixel_index2 <= 620)) || pixel_index2 == 631 || ((pixel_index2 >= 637) && (pixel_index2 <= 640)) || ((pixel_index2 >= 645) && (pixel_index2 <= 646)) || pixel_index2 == 651 || pixel_index2 == 657 || pixel_index2 == 670 || ((pixel_index2 >= 672) && (pixel_index2 <= 673)) || pixel_index2 == 676 || ((pixel_index2 >= 678) && (pixel_index2 <= 679)) || pixel_index2 == 691 || pixel_index2 == 694 || pixel_index2 == 696 || pixel_index2 == 700 || pixel_index2 == 704 || pixel_index2 == 707 || ((pixel_index2 >= 715) && (pixel_index2 <= 716)) || ((pixel_index2 >= 726) && (pixel_index2 <= 727)) || ((pixel_index2 >= 733) && (pixel_index2 <= 736)) || ((pixel_index2 >= 741) && (pixel_index2 <= 742)) || pixel_index2 == 744 || pixel_index2 == 766 || pixel_index2 == 769 || ((pixel_index2 >= 774) && (pixel_index2 <= 775)) || pixel_index2 == 779 || pixel_index2 == 783 || pixel_index2 == 787 || pixel_index2 == 790 || pixel_index2 == 800 || pixel_index2 == 803 || pixel_index2 == 811 || pixel_index2 == 822 || pixel_index2 == 825 || ((pixel_index2 >= 829) && (pixel_index2 <= 831)) || pixel_index2 == 841 || ((pixel_index2 >= 844) && (pixel_index2 <= 846)) || pixel_index2 == 853 || pixel_index2 == 862 || pixel_index2 == 865 || pixel_index2 == 871 || pixel_index2 == 879 || pixel_index2 == 883 || pixel_index2 == 896 || pixel_index2 == 899 || pixel_index2 == 918 || pixel_index2 == 921 || ((pixel_index2 >= 925) && (pixel_index2 <= 927)) || pixel_index2 == 937 || pixel_index2 == 940 || pixel_index2 == 955 || pixel_index2 == 958 || pixel_index2 == 961 || pixel_index2 == 965 || pixel_index2 == 967 || ((pixel_index2 >= 970) && (pixel_index2 <= 971)) || pixel_index2 == 975 || pixel_index2 == 979 || pixel_index2 == 982 || pixel_index2 == 998 || ((pixel_index2 >= 1002) && (pixel_index2 <= 1003)) || pixel_index2 == 1014 || ((pixel_index2 >= 1020) && (pixel_index2 <= 1023)) || ((pixel_index2 >= 1041) && (pixel_index2 <= 1042)) || pixel_index2 == 1054 || pixel_index2 == 1061 || ((pixel_index2 >= 1064) && (pixel_index2 <= 1065)) || ((pixel_index2 >= 1068) && (pixel_index2 <= 1072)) || ((pixel_index2 >= 1074) && (pixel_index2 <= 1075)) || ((pixel_index2 >= 1078) && (pixel_index2 <= 1082)) || ((pixel_index2 >= 1093) && (pixel_index2 <= 1095)) || pixel_index2 == 1097 || pixel_index2 == 1100 || pixel_index2 == 1103 || pixel_index2 == 1111 || ((pixel_index2 >= 1113) && (pixel_index2 <= 1114)) || ((pixel_index2 >= 1116) && (pixel_index2 <= 1120)) || ((pixel_index2 >= 1122) && (pixel_index2 <= 1123)) || ((pixel_index2 >= 1125) && (pixel_index2 <= 1126)) || ((pixel_index2 >= 1128) && (pixel_index2 <= 1132)) || ((pixel_index2 >= 1137) && (pixel_index2 <= 1138)) || pixel_index2 == 1144 || pixel_index2 == 1156 || ((pixel_index2 >= 1199) && (pixel_index2 <= 1242)) || pixel_index2 == 1252 || ((pixel_index2 >= 1296) && (pixel_index2 <= 1306)) || ((pixel_index2 >= 1311) && (pixel_index2 <= 1333)) || ((pixel_index2 >= 1335) && (pixel_index2 <= 1338)) || pixel_index2 == 1349 || ((pixel_index2 >= 1394) && (pixel_index2 <= 1403)) || ((pixel_index2 >= 1408) && (pixel_index2 <= 1429)) || ((pixel_index2 >= 1431) && (pixel_index2 <= 1434)) || pixel_index2 == 1445 || ((pixel_index2 >= 1493) && (pixel_index2 <= 1501)) || pixel_index2 == 1505 || ((pixel_index2 >= 1513) && (pixel_index2 <= 1531)) || ((pixel_index2 >= 1536) && (pixel_index2 <= 1538)) || pixel_index2 == 1541 || ((pixel_index2 >= 1592) && (pixel_index2 <= 1598)) || ((pixel_index2 >= 1610) && (pixel_index2 <= 1627)) || ((pixel_index2 >= 1632) && (pixel_index2 <= 1633)) || pixel_index2 == 1637 || ((pixel_index2 >= 1689) && (pixel_index2 <= 1694)) || ((pixel_index2 >= 1706) && (pixel_index2 <= 1724)) || pixel_index2 == 1728 || pixel_index2 == 1733 || ((pixel_index2 >= 1785) && (pixel_index2 <= 1791)) || ((pixel_index2 >= 1804) && (pixel_index2 <= 1815)) || ((pixel_index2 >= 1817) && (pixel_index2 <= 1820)) || pixel_index2 == 1829 || ((pixel_index2 >= 1881) && (pixel_index2 <= 1886)) || ((pixel_index2 >= 1900) && (pixel_index2 <= 1916)) || pixel_index2 == 1925 || ((pixel_index2 >= 1977) && (pixel_index2 <= 1982)) || ((pixel_index2 >= 1996) && (pixel_index2 <= 2008)) || ((pixel_index2 >= 2011) && (pixel_index2 <= 2012)) || pixel_index2 == 2020 || ((pixel_index2 >= 2073) && (pixel_index2 <= 2078)) || ((pixel_index2 >= 2093) && (pixel_index2 <= 2103)) || ((pixel_index2 >= 2107) && (pixel_index2 <= 2109)) || pixel_index2 == 2116 || ((pixel_index2 >= 2169) && (pixel_index2 <= 2173)) || ((pixel_index2 >= 2191) && (pixel_index2 <= 2198)) || ((pixel_index2 >= 2204) && (pixel_index2 <= 2205)) || pixel_index2 == 2212 || ((pixel_index2 >= 2266) && (pixel_index2 <= 2269)) || ((pixel_index2 >= 2290) && (pixel_index2 <= 2294)) || ((pixel_index2 >= 2300) && (pixel_index2 <= 2301)) || ((pixel_index2 >= 2387) && (pixel_index2 <= 2389)) || pixel_index2 == 2397 || ((pixel_index2 >= 2484) && (pixel_index2 <= 2485)) || ((pixel_index2 >= 2493) && (pixel_index2 <= 2494)) || pixel_index2 == 2499 || ((pixel_index2 >= 2589) && (pixel_index2 <= 2590)) || pixel_index2 == 2595 || ((pixel_index2 >= 2685) && (pixel_index2 <= 2686)) || ((pixel_index2 >= 2688) && (pixel_index2 <= 2691)) || ((pixel_index2 >= 2781) && (pixel_index2 <= 2782)) || ((pixel_index2 >= 2784) && (pixel_index2 <= 2785)) || pixel_index2 == 2787 || pixel_index2 == 2867 || pixel_index2 == 2878 || ((pixel_index2 >= 2901) && (pixel_index2 <= 2910)) || ((pixel_index2 >= 2944) && (pixel_index2 <= 2948)) || pixel_index2 == 2963 || pixel_index2 == 2974 || pixel_index2 == 2976 || ((pixel_index2 >= 2995) && (pixel_index2 <= 2999)) || ((pixel_index2 >= 3006) && (pixel_index2 <= 3008)) || ((pixel_index2 >= 3040) && (pixel_index2 <= 3058)) || pixel_index2 == 3070 || pixel_index2 == 3074 || ((pixel_index2 >= 3090) && (pixel_index2 <= 3093)) || ((pixel_index2 >= 3104) && (pixel_index2 <= 3105)) || ((pixel_index2 >= 3137) && (pixel_index2 <= 3154)) || pixel_index2 == 3166 || pixel_index2 == 3170 || ((pixel_index2 >= 3186) && (pixel_index2 <= 3188)) || ((pixel_index2 >= 3200) && (pixel_index2 <= 3201)) || ((pixel_index2 >= 3232) && (pixel_index2 <= 3239)) || ((pixel_index2 >= 3246) && (pixel_index2 <= 3250)) || pixel_index2 == 3262 || ((pixel_index2 >= 3282) && (pixel_index2 <= 3284)) || ((pixel_index2 >= 3297) && (pixel_index2 <= 3298)) || ((pixel_index2 >= 3328) && (pixel_index2 <= 3331)) || ((pixel_index2 >= 3344) && (pixel_index2 <= 3347)) || pixel_index2 == 3358 || ((pixel_index2 >= 3378) && (pixel_index2 <= 3380)) || ((pixel_index2 >= 3393) && (pixel_index2 <= 3394)) || ((pixel_index2 >= 3424) && (pixel_index2 <= 3427)) || ((pixel_index2 >= 3441) && (pixel_index2 <= 3443)) || pixel_index2 == 3454 || ((pixel_index2 >= 3474) && (pixel_index2 <= 3477)) || ((pixel_index2 >= 3489) && (pixel_index2 <= 3490)) || ((pixel_index2 >= 3521) && (pixel_index2 <= 3523)) || ((pixel_index2 >= 3537) && (pixel_index2 <= 3540)) || pixel_index2 == 3550 || ((pixel_index2 >= 3570) && (pixel_index2 <= 3573)) || ((pixel_index2 >= 3584) && (pixel_index2 <= 3585)) || ((pixel_index2 >= 3618) && (pixel_index2 <= 3619)) || ((pixel_index2 >= 3633) && (pixel_index2 <= 3637)) || pixel_index2 == 3646 || ((pixel_index2 >= 3666) && (pixel_index2 <= 3669)) || ((pixel_index2 >= 3678) && (pixel_index2 <= 3680)) || ((pixel_index2 >= 3715) && (pixel_index2 <= 3717)) || ((pixel_index2 >= 3729) && (pixel_index2 <= 3733)) || pixel_index2 == 3742 || pixel_index2 == 3746 || ((pixel_index2 >= 3765) && (pixel_index2 <= 3773)) || ((pixel_index2 >= 3812) && (pixel_index2 <= 3815)) || ((pixel_index2 >= 3825) && (pixel_index2 <= 3829)) || pixel_index2 == 3838 || pixel_index2 == 3842 || ((pixel_index2 >= 3910) && (pixel_index2 <= 3913)) || ((pixel_index2 >= 3919) && (pixel_index2 <= 3925)) || pixel_index2 == 3934 || pixel_index2 == 3938 || ((pixel_index2 >= 4008) && (pixel_index2 <= 4018)) || ((pixel_index2 >= 4029) && (pixel_index2 <= 4030)) || pixel_index2 == 4034 || pixel_index2 == 4125 || pixel_index2 == 4130 || pixel_index2 == 4221 || pixel_index2 == 4226 || pixel_index2 == 4316 || pixel_index2 == 4322 || pixel_index2 == 4412 || pixel_index2 == 4418 || pixel_index2 == 4509 || pixel_index2 == 4513 || pixel_index2 == 4606 || pixel_index2 == 4609 || pixel_index2 == 4699 || pixel_index2 == 4702 || pixel_index2 == 4705 || ((pixel_index2 >= 4793) && (pixel_index2 <= 4795)) || pixel_index2 == 4798 || pixel_index2 == 4801 || ((pixel_index2 >= 4885) && (pixel_index2 <= 4891)) || pixel_index2 == 4894 || pixel_index2 == 4897 || ((pixel_index2 >= 4920) && (pixel_index2 <= 4923)) || pixel_index2 == 4925 || pixel_index2 == 4927 || pixel_index2 == 4929 || ((pixel_index2 >= 4933) && (pixel_index2 <= 4936)) || pixel_index2 == 4940 || pixel_index2 == 4945 || ((pixel_index2 >= 4949) && (pixel_index2 <= 4953)) || pixel_index2 == 4955 || pixel_index2 == 4958 || pixel_index2 == 4961 || pixel_index2 == 4963 || pixel_index2 == 4968 || ((pixel_index2 >= 4978) && (pixel_index2 <= 4986)) || pixel_index2 == 4990 || pixel_index2 == 4993 || pixel_index2 == 5016 || pixel_index2 == 5024 || ((pixel_index2 >= 5027) && (pixel_index2 <= 5028)) || ((pixel_index2 >= 5034) && (pixel_index2 <= 5035)) || pixel_index2 == 5044 || ((pixel_index2 >= 5050) && (pixel_index2 <= 5051)) || ((pixel_index2 >= 5074) && (pixel_index2 <= 5081)) || pixel_index2 == 5086 || pixel_index2 == 5089 || pixel_index2 == 5112 || pixel_index2 == 5120 || pixel_index2 == 5123 || pixel_index2 == 5127 || pixel_index2 == 5130 || pixel_index2 == 5134 || pixel_index2 == 5143 || ((pixel_index2 >= 5146) && (pixel_index2 <= 5147)) || pixel_index2 == 5154 || pixel_index2 == 5157 || ((pixel_index2 >= 5170) && (pixel_index2 <= 5174)) || pixel_index2 == 5183 || pixel_index2 == 5186 || pixel_index2 == 5208 || pixel_index2 == 5216 || pixel_index2 == 5219 || pixel_index2 == 5223 || pixel_index2 == 5226 || pixel_index2 == 5236 || pixel_index2 == 5239 || pixel_index2 == 5243 || pixel_index2 == 5250 || ((pixel_index2 >= 5267) && (pixel_index2 <= 5270)) || pixel_index2 == 5279 || pixel_index2 == 5282 || pixel_index2 == 5304 || pixel_index2 == 5315 || pixel_index2 == 5319 || pixel_index2 == 5322 || pixel_index2 == 5332 || pixel_index2 == 5335 || pixel_index2 == 5339 || pixel_index2 == 5346 || pixel_index2 == 5375 || pixel_index2 == 5377 || pixel_index2 == 5400 || pixel_index2 == 5411 || pixel_index2 == 5415 || pixel_index2 == 5418 || pixel_index2 == 5428 || pixel_index2 == 5431 || pixel_index2 == 5435 || pixel_index2 == 5442 || ((pixel_index2 >= 5471) && (pixel_index2 <= 5473)) || pixel_index2 == 5496 || pixel_index2 == 5507 || pixel_index2 == 5511 || pixel_index2 == 5514 || pixel_index2 == 5524 || pixel_index2 == 5527 || pixel_index2 == 5531 || pixel_index2 == 5538 || ((pixel_index2 >= 5582) && (pixel_index2 <= 5584)) || ((pixel_index2 >= 5589) && (pixel_index2 <= 5591)) || pixel_index2 == 5603 || pixel_index2 == 5607 || pixel_index2 == 5610 || pixel_index2 == 5620 || pixel_index2 == 5623 || pixel_index2 == 5627 || pixel_index2 == 5634 || ((pixel_index2 >= 5674) && (pixel_index2 <= 5678)) || pixel_index2 == 5688 || pixel_index2 == 5699 || pixel_index2 == 5703 || pixel_index2 == 5706 || pixel_index2 == 5716 || pixel_index2 == 5719 || pixel_index2 == 5723 || pixel_index2 == 5730 || pixel_index2 == 5737 || ((pixel_index2 >= 5741) && (pixel_index2 <= 5746)) || ((pixel_index2 >= 5768) && (pixel_index2 <= 5770)) || pixel_index2 == 5792 || ((pixel_index2 >= 5795) && (pixel_index2 <= 5796)) || pixel_index2 == 5803 || pixel_index2 == 5811 || pixel_index2 == 5818 || pixel_index2 == 5832 || ((pixel_index2 >= 5837) && (pixel_index2 <= 5843)) || ((pixel_index2 >= 5862) && (pixel_index2 <= 5865)) || pixel_index2 == 5891 || pixel_index2 == 5893 || pixel_index2 == 5897 || pixel_index2 == 5900 || pixel_index2 == 5909 || pixel_index2 == 5913 || pixel_index2 == 5916 || pixel_index2 == 5921 || pixel_index2 == 5923 || pixel_index2 == 5928 || ((pixel_index2 >= 5932) && (pixel_index2 <= 5944)) || ((pixel_index2 >= 5956) && (pixel_index2 <= 5958)) || ((pixel_index2 >= 6028) && (pixel_index2 <= 6043)) || ((pixel_index2 >= 6051) && (pixel_index2 <= 6053)) || ((pixel_index2 >= 6071) && (pixel_index2 <= 6072)) || (pixel_index2 >= 6124) && (pixel_index2 <= 6141)) oled_data2 = 16'b0101001010001010;
        else if (((pixel_index2 >= 29) && (pixel_index2 <= 31)) || pixel_index2 == 99 || ((pixel_index2 >= 104) && (pixel_index2 <= 105)) || pixel_index2 == 114 || pixel_index2 == 124 || pixel_index2 == 126 || pixel_index2 == 152 || pixel_index2 == 170 || pixel_index2 == 204 || ((pixel_index2 >= 222) && (pixel_index2 <= 223)) || pixel_index2 == 230 || ((pixel_index2 >= 318) && (pixel_index2 <= 319)) || pixel_index2 == 420 || pixel_index2 == 453 || pixel_index2 == 480 || pixel_index2 == 516 || pixel_index2 == 612 || pixel_index2 == 708 || pixel_index2 == 749 || pixel_index2 == 778 || pixel_index2 == 804 || pixel_index2 == 922 || pixel_index2 == 993 || pixel_index2 == 1015 || pixel_index2 == 1089 || ((pixel_index2 >= 1171) && (pixel_index2 <= 1172)) || pixel_index2 == 1194 || ((pixel_index2 >= 1265) && (pixel_index2 <= 1269)) || pixel_index2 == 1350 || ((pixel_index2 >= 1361) && (pixel_index2 <= 1365)) || pixel_index2 == 1387 || pixel_index2 == 1446 || ((pixel_index2 >= 1456) && (pixel_index2 <= 1461)) || pixel_index2 == 1483 || pixel_index2 == 1542 || ((pixel_index2 >= 1552) && (pixel_index2 <= 1557)) || ((pixel_index2 >= 1579) && (pixel_index2 <= 1581)) || pixel_index2 == 1638 || ((pixel_index2 >= 1648) && (pixel_index2 <= 1653)) || pixel_index2 == 1677 || pixel_index2 == 1734 || ((pixel_index2 >= 1744) && (pixel_index2 <= 1749)) || ((pixel_index2 >= 1774) && (pixel_index2 <= 1775)) || ((pixel_index2 >= 1840) && (pixel_index2 <= 1845)) || ((pixel_index2 >= 1871) && (pixel_index2 <= 1872)) || ((pixel_index2 >= 1890) && (pixel_index2 <= 1896)) || ((pixel_index2 >= 1936) && (pixel_index2 <= 1941)) || ((pixel_index2 >= 1968) && (pixel_index2 <= 1969)) || ((pixel_index2 >= 1985) && (pixel_index2 <= 1986)) || ((pixel_index2 >= 1988) && (pixel_index2 <= 1993)) || ((pixel_index2 >= 2032) && (pixel_index2 <= 2037)) || ((pixel_index2 >= 2066) && (pixel_index2 <= 2067)) || ((pixel_index2 >= 2081) && (pixel_index2 <= 2083)) || ((pixel_index2 >= 2085) && (pixel_index2 <= 2091)) || pixel_index2 == 2117 || ((pixel_index2 >= 2128) && (pixel_index2 <= 2133)) || ((pixel_index2 >= 2163) && (pixel_index2 <= 2164)) || pixel_index2 == 2178 || ((pixel_index2 >= 2186) && (pixel_index2 <= 2188)) || pixel_index2 == 2213 || ((pixel_index2 >= 2224) && (pixel_index2 <= 2230)) || pixel_index2 == 2260 || pixel_index2 == 2272 || ((pixel_index2 >= 2284) && (pixel_index2 <= 2286)) || ((pixel_index2 >= 2320) && (pixel_index2 <= 2326)) || pixel_index2 == 2368 || ((pixel_index2 >= 2381) && (pixel_index2 <= 2383)) || ((pixel_index2 >= 2416) && (pixel_index2 <= 2423)) || pixel_index2 == 2454 || pixel_index2 == 2464 || ((pixel_index2 >= 2478) && (pixel_index2 <= 2480)) || pixel_index2 == 2500 || ((pixel_index2 >= 2511) && (pixel_index2 <= 2519)) || ((pixel_index2 >= 2550) && (pixel_index2 <= 2551)) || pixel_index2 == 2560 || ((pixel_index2 >= 2575) && (pixel_index2 <= 2577)) || pixel_index2 == 2596 || ((pixel_index2 >= 2607) && (pixel_index2 <= 2615)) || pixel_index2 == 2648 || ((pixel_index2 >= 2655) && (pixel_index2 <= 2657)) || ((pixel_index2 >= 2672) && (pixel_index2 <= 2673)) || ((pixel_index2 >= 2703) && (pixel_index2 <= 2711)) || ((pixel_index2 >= 2743) && (pixel_index2 <= 2744)) || ((pixel_index2 >= 2751) && (pixel_index2 <= 2757)) || ((pixel_index2 >= 2767) && (pixel_index2 <= 2769)) || ((pixel_index2 >= 2799) && (pixel_index2 <= 2802)) || ((pixel_index2 >= 2804) && (pixel_index2 <= 2808)) || ((pixel_index2 >= 2813) && (pixel_index2 <= 2815)) || ((pixel_index2 >= 2838) && (pixel_index2 <= 2847)) || ((pixel_index2 >= 2855) && (pixel_index2 <= 2857)) || ((pixel_index2 >= 2863) && (pixel_index2 <= 2864)) || ((pixel_index2 >= 2895) && (pixel_index2 <= 2897)) || pixel_index2 == 2914 || ((pixel_index2 >= 2934) && (pixel_index2 <= 2941)) || ((pixel_index2 >= 2956) && (pixel_index2 <= 2959)) || ((pixel_index2 >= 2991) && (pixel_index2 <= 2993)) || pixel_index2 == 3011 || ((pixel_index2 >= 3030) && (pixel_index2 <= 3037)) || pixel_index2 == 3075 || ((pixel_index2 >= 3088) && (pixel_index2 <= 3089)) || pixel_index2 == 3108 || ((pixel_index2 >= 3127) && (pixel_index2 <= 3133)) || pixel_index2 == 3184 || ((pixel_index2 >= 3223) && (pixel_index2 <= 3229)) || pixel_index2 == 3280 || ((pixel_index2 >= 3319) && (pixel_index2 <= 3325)) || ((pixel_index2 >= 3349) && (pixel_index2 <= 3350)) || pixel_index2 == 3376 || pixel_index2 == 3397 || ((pixel_index2 >= 3416) && (pixel_index2 <= 3421)) || ((pixel_index2 >= 3446) && (pixel_index2 <= 3447)) || pixel_index2 == 3472 || ((pixel_index2 >= 3493) && (pixel_index2 <= 3494)) || ((pixel_index2 >= 3512) && (pixel_index2 <= 3518)) || ((pixel_index2 >= 3543) && (pixel_index2 <= 3544)) || ((pixel_index2 >= 3590) && (pixel_index2 <= 3591)) || ((pixel_index2 >= 3608) && (pixel_index2 <= 3613)) || pixel_index2 == 3665 || ((pixel_index2 >= 3685) && (pixel_index2 <= 3689)) || ((pixel_index2 >= 3705) && (pixel_index2 <= 3709)) || ((pixel_index2 >= 3736) && (pixel_index2 <= 3740)) || pixel_index2 == 3747 || pixel_index2 == 3777 || ((pixel_index2 >= 3780) && (pixel_index2 <= 3787)) || ((pixel_index2 >= 3802) && (pixel_index2 <= 3806)) || ((pixel_index2 >= 3831) && (pixel_index2 <= 3836)) || pixel_index2 == 3843 || ((pixel_index2 >= 3862) && (pixel_index2 <= 3871)) || ((pixel_index2 >= 3873) && (pixel_index2 <= 3884)) || ((pixel_index2 >= 3898) && (pixel_index2 <= 3904)) || ((pixel_index2 >= 3927) && (pixel_index2 <= 3932)) || pixel_index2 == 3940 || ((pixel_index2 >= 3964) && (pixel_index2 <= 3981)) || ((pixel_index2 >= 3996) && (pixel_index2 <= 4001)) || ((pixel_index2 >= 4022) && (pixel_index2 <= 4028)) || pixel_index2 == 4036 || ((pixel_index2 >= 4060) && (pixel_index2 <= 4078)) || ((pixel_index2 >= 4095) && (pixel_index2 <= 4099)) || ((pixel_index2 >= 4118) && (pixel_index2 <= 4124)) || ((pixel_index2 >= 4132) && (pixel_index2 <= 4133)) || ((pixel_index2 >= 4157) && (pixel_index2 <= 4175)) || ((pixel_index2 >= 4192) && (pixel_index2 <= 4195)) || ((pixel_index2 >= 4214) && (pixel_index2 <= 4219)) || ((pixel_index2 >= 4229) && (pixel_index2 <= 4230)) || ((pixel_index2 >= 4253) && (pixel_index2 <= 4258)) || ((pixel_index2 >= 4261) && (pixel_index2 <= 4272)) || ((pixel_index2 >= 4289) && (pixel_index2 <= 4292)) || pixel_index2 == 4301 || ((pixel_index2 >= 4310) && (pixel_index2 <= 4315)) || ((pixel_index2 >= 4325) && (pixel_index2 <= 4329)) || ((pixel_index2 >= 4359) && (pixel_index2 <= 4369)) || ((pixel_index2 >= 4384) && (pixel_index2 <= 4397)) || ((pixel_index2 >= 4405) && (pixel_index2 <= 4411)) || ((pixel_index2 >= 4420) && (pixel_index2 <= 4425)) || ((pixel_index2 >= 4456) && (pixel_index2 <= 4465)) || ((pixel_index2 >= 4478) && (pixel_index2 <= 4494)) || ((pixel_index2 >= 4500) && (pixel_index2 <= 4503)) || pixel_index2 == 4505 || ((pixel_index2 >= 4516) && (pixel_index2 <= 4519)) || ((pixel_index2 >= 4521) && (pixel_index2 <= 4522)) || pixel_index2 == 4551 || ((pixel_index2 >= 4553) && (pixel_index2 <= 4561)) || ((pixel_index2 >= 4568) && (pixel_index2 <= 4591)) || ((pixel_index2 >= 4596) && (pixel_index2 <= 4598)) || ((pixel_index2 >= 4611) && (pixel_index2 <= 4615)) || ((pixel_index2 >= 4618) && (pixel_index2 <= 4620)) || ((pixel_index2 >= 4647) && (pixel_index2 <= 4658)) || ((pixel_index2 >= 4664) && (pixel_index2 <= 4687)) || ((pixel_index2 >= 4693) && (pixel_index2 <= 4694)) || ((pixel_index2 >= 4707) && (pixel_index2 <= 4711)) || ((pixel_index2 >= 4716) && (pixel_index2 <= 4718)) || ((pixel_index2 >= 4745) && (pixel_index2 <= 4749)) || ((pixel_index2 >= 4753) && (pixel_index2 <= 4754)) || ((pixel_index2 >= 4760) && (pixel_index2 <= 4784)) || ((pixel_index2 >= 4803) && (pixel_index2 <= 4808)) || ((pixel_index2 >= 4812) && (pixel_index2 <= 4817)) || pixel_index2 == 4851 || ((pixel_index2 >= 4855) && (pixel_index2 <= 4868)) || ((pixel_index2 >= 4872) && (pixel_index2 <= 4879)) || ((pixel_index2 >= 4899) && (pixel_index2 <= 4906)) || ((pixel_index2 >= 4911) && (pixel_index2 <= 4915)) || pixel_index2 == 4939 || pixel_index2 == 4954 || pixel_index2 == 4962 || ((pixel_index2 >= 4969) && (pixel_index2 <= 4974)) || ((pixel_index2 >= 4996) && (pixel_index2 <= 5000)) || ((pixel_index2 >= 5010) && (pixel_index2 <= 5012)) || ((pixel_index2 >= 5064) && (pixel_index2 <= 5069)) || ((pixel_index2 >= 5092) && (pixel_index2 <= 5096)) || ((pixel_index2 >= 5106) && (pixel_index2 <= 5108)) || ((pixel_index2 >= 5160) && (pixel_index2 <= 5165)) || ((pixel_index2 >= 5188) && (pixel_index2 <= 5192)) || ((pixel_index2 >= 5202) && (pixel_index2 <= 5204)) || pixel_index2 == 5256 || ((pixel_index2 >= 5258) && (pixel_index2 <= 5260)) || ((pixel_index2 >= 5284) && (pixel_index2 <= 5288)) || ((pixel_index2 >= 5297) && (pixel_index2 <= 5299)) || pixel_index2 == 5352 || ((pixel_index2 >= 5355) && (pixel_index2 <= 5360)) || pixel_index2 == 5362 || ((pixel_index2 >= 5379) && (pixel_index2 <= 5383)) || ((pixel_index2 >= 5393) && (pixel_index2 <= 5395)) || pixel_index2 == 5448 || ((pixel_index2 >= 5456) && (pixel_index2 <= 5464)) || ((pixel_index2 >= 5475) && (pixel_index2 <= 5478)) || ((pixel_index2 >= 5491) && (pixel_index2 <= 5492)) || pixel_index2 == 5544 || ((pixel_index2 >= 5553) && (pixel_index2 <= 5560)) || ((pixel_index2 >= 5569) && (pixel_index2 <= 5572)) || pixel_index2 == 5596 || pixel_index2 == 5640 || ((pixel_index2 >= 5646) && (pixel_index2 <= 5660)) || pixel_index2 == 5662 || ((pixel_index2 >= 5664) && (pixel_index2 <= 5668)) || pixel_index2 == 5722 || pixel_index2 == 5738 || ((pixel_index2 >= 5748) && (pixel_index2 <= 5758)) || ((pixel_index2 >= 5760) && (pixel_index2 <= 5763)) || ((pixel_index2 >= 5846) && (pixel_index2 <= 5854)) || ((pixel_index2 >= 5856) && (pixel_index2 <= 5858)) || ((pixel_index2 >= 5947) && (pixel_index2 <= 5950)) || ((pixel_index2 >= 5952) && (pixel_index2 <= 5953)) || ((pixel_index2 >= 6045) && (pixel_index2 <= 6046)) || (pixel_index2 >= 6048) && (pixel_index2 <= 6049)) oled_data2 = 16'b1010010100001010;
        else if (pixel_index2 == 149 || pixel_index2 == 220 || pixel_index2 == 246 || pixel_index2 == 280 || pixel_index2 == 283 || pixel_index2 == 287 || pixel_index2 == 376 || pixel_index2 == 383 || pixel_index2 == 472 || pixel_index2 == 479 || pixel_index2 == 512 || pixel_index2 == 575 || pixel_index2 == 608 || pixel_index2 == 630 || pixel_index2 == 636 || pixel_index2 == 767 || ((pixel_index2 >= 863) && (pixel_index2 <= 864)) || pixel_index2 == 886 || ((pixel_index2 >= 959) && (pixel_index2 <= 960)) || pixel_index2 == 988 || pixel_index2 == 1007 || ((pixel_index2 >= 1055) && (pixel_index2 <= 1056)) || pixel_index2 == 1060 || ((pixel_index2 >= 1101) && (pixel_index2 <= 1102)) || ((pixel_index2 >= 1104) && (pixel_index2 <= 1110)) || ((pixel_index2 >= 1140) && (pixel_index2 <= 1141)) || pixel_index2 == 1145 || ((pixel_index2 >= 1151) && (pixel_index2 <= 1154)) || ((pixel_index2 >= 1247) && (pixel_index2 <= 1250)) || pixel_index2 == 1343 || pixel_index2 == 1439 || pixel_index2 == 1535 || pixel_index2 == 1631 || ((pixel_index2 >= 1726) && (pixel_index2 <= 1727)) || pixel_index2 == 1730 || ((pixel_index2 >= 1826) && (pixel_index2 <= 1827)) || ((pixel_index2 >= 1920) && (pixel_index2 <= 1923)) || ((pixel_index2 >= 2015) && (pixel_index2 <= 2019)) || ((pixel_index2 >= 2111) && (pixel_index2 <= 2115)) || ((pixel_index2 >= 2207) && (pixel_index2 <= 2211)) || ((pixel_index2 >= 2303) && (pixel_index2 <= 2306)) || ((pixel_index2 >= 2399) && (pixel_index2 <= 2402)) || ((pixel_index2 >= 2495) && (pixel_index2 <= 2497)) || pixel_index2 == 2591 || pixel_index2 == 2687 || pixel_index2 == 3002 || ((pixel_index2 >= 3096) && (pixel_index2 <= 3102)) || pixel_index2 == 3168 || pixel_index2 == 3190 || pixel_index2 == 3192 || ((pixel_index2 >= 3197) && (pixel_index2 <= 3198)) || pixel_index2 == 3244 || ((pixel_index2 >= 3264) && (pixel_index2 <= 3265)) || pixel_index2 == 3285 || ((pixel_index2 >= 3293) && (pixel_index2 <= 3295)) || ((pixel_index2 >= 3333) && (pixel_index2 <= 3335)) || pixel_index2 == 3343 || ((pixel_index2 >= 3360) && (pixel_index2 <= 3361)) || pixel_index2 == 3381 || ((pixel_index2 >= 3383) && (pixel_index2 <= 3386)) || ((pixel_index2 >= 3389) && (pixel_index2 <= 3391)) || ((pixel_index2 >= 3428) && (pixel_index2 <= 3430)) || pixel_index2 == 3439 || ((pixel_index2 >= 3456) && (pixel_index2 <= 3457)) || ((pixel_index2 >= 3478) && (pixel_index2 <= 3480)) || pixel_index2 == 3482 || ((pixel_index2 >= 3485) && (pixel_index2 <= 3487)) || ((pixel_index2 >= 3524) && (pixel_index2 <= 3526)) || ((pixel_index2 >= 3552) && (pixel_index2 <= 3553)) || ((pixel_index2 >= 3574) && (pixel_index2 <= 3575)) || ((pixel_index2 >= 3578) && (pixel_index2 <= 3579)) || ((pixel_index2 >= 3581) && (pixel_index2 <= 3582)) || ((pixel_index2 >= 3621) && (pixel_index2 <= 3623)) || ((pixel_index2 >= 3625) && (pixel_index2 <= 3626)) || ((pixel_index2 >= 3648) && (pixel_index2 <= 3649)) || ((pixel_index2 >= 3670) && (pixel_index2 <= 3676)) || ((pixel_index2 >= 3719) && (pixel_index2 <= 3723)) || pixel_index2 == 3728 || ((pixel_index2 >= 3743) && (pixel_index2 <= 3745)) || ((pixel_index2 >= 3817) && (pixel_index2 <= 3824)) || ((pixel_index2 >= 3839) && (pixel_index2 <= 3841)) || pixel_index2 == 3936 || pixel_index2 == 4032 || pixel_index2 == 4126 || pixel_index2 == 4128 || pixel_index2 == 4224 || pixel_index2 == 4320 || pixel_index2 == 4416 || pixel_index2 == 4510 || pixel_index2 == 4512 || ((pixel_index2 >= 4607) && (pixel_index2 <= 4608)) || pixel_index2 == 4704 || pixel_index2 == 4800 || pixel_index2 == 4896 || ((pixel_index2 >= 4941) && (pixel_index2 <= 4944)) || pixel_index2 == 4960 || ((pixel_index2 >= 4964) && (pixel_index2 <= 4967)) || pixel_index2 == 4992 || pixel_index2 == 5019 || pixel_index2 == 5088 || pixel_index2 == 5140 || pixel_index2 == 5185 || pixel_index2 == 5280 || pixel_index2 == 5586 || pixel_index2 == 5680 || ((pixel_index2 >= 5684) && (pixel_index2 <= 5685)) || pixel_index2 == 5772 || ((pixel_index2 >= 5774) && (pixel_index2 <= 5776)) || pixel_index2 == 5834 || pixel_index2 == 5867 || pixel_index2 == 5964 || ((pixel_index2 >= 6054) && (pixel_index2 <= 6056)) || (pixel_index2 >= 6082) && (pixel_index2 <= 6085)) oled_data2 = 16'b0101000000000000;
        else if (pixel_index2 == 156 || pixel_index2 == 177 || pixel_index2 == 202 || pixel_index2 == 298 || pixel_index2 == 394 || pixel_index2 == 540 || pixel_index2 == 561 || pixel_index2 == 569 || pixel_index2 == 652 || pixel_index2 == 658 || pixel_index2 == 671 || pixel_index2 == 682 || pixel_index2 == 743 || pixel_index2 == 753 || pixel_index2 == 768 || pixel_index2 == 908 || pixel_index2 == 999 || pixel_index2 == 1073 || ((pixel_index2 >= 1076) && (pixel_index2 <= 1077)) || pixel_index2 == 1083 || pixel_index2 == 1090 || pixel_index2 == 1096 || pixel_index2 == 1121 || ((pixel_index2 >= 1133) && (pixel_index2 <= 1136)) || ((pixel_index2 >= 1142) && (pixel_index2 <= 1143)) || pixel_index2 == 1155 || ((pixel_index2 >= 1243) && (pixel_index2 <= 1246)) || pixel_index2 == 1251 || ((pixel_index2 >= 1339) && (pixel_index2 <= 1342)) || ((pixel_index2 >= 1344) && (pixel_index2 <= 1348)) || ((pixel_index2 >= 1435) && (pixel_index2 <= 1438)) || ((pixel_index2 >= 1440) && (pixel_index2 <= 1444)) || ((pixel_index2 >= 1532) && (pixel_index2 <= 1534)) || ((pixel_index2 >= 1539) && (pixel_index2 <= 1540)) || ((pixel_index2 >= 1628) && (pixel_index2 <= 1630)) || ((pixel_index2 >= 1634) && (pixel_index2 <= 1636)) || pixel_index2 == 1725 || pixel_index2 == 1729 || ((pixel_index2 >= 1731) && (pixel_index2 <= 1732)) || ((pixel_index2 >= 1821) && (pixel_index2 <= 1822)) || ((pixel_index2 >= 1824) && (pixel_index2 <= 1825)) || pixel_index2 == 1828 || ((pixel_index2 >= 1917) && (pixel_index2 <= 1918)) || pixel_index2 == 1924 || ((pixel_index2 >= 2013) && (pixel_index2 <= 2014)) || pixel_index2 == 2110 || pixel_index2 == 2206 || pixel_index2 == 2302 || pixel_index2 == 2307 || pixel_index2 == 2398 || pixel_index2 == 2403 || pixel_index2 == 2498 || ((pixel_index2 >= 2592) && (pixel_index2 <= 2594)) || pixel_index2 == 2783 || pixel_index2 == 2786 || ((pixel_index2 >= 2879) && (pixel_index2 <= 2882)) || pixel_index2 == 2975 || ((pixel_index2 >= 2977) && (pixel_index2 <= 2978)) || ((pixel_index2 >= 3000) && (pixel_index2 <= 3001)) || ((pixel_index2 >= 3003) && (pixel_index2 <= 3005)) || ((pixel_index2 >= 3071) && (pixel_index2 <= 3073)) || ((pixel_index2 >= 3094) && (pixel_index2 <= 3095)) || pixel_index2 == 3103 || pixel_index2 == 3167 || pixel_index2 == 3169 || pixel_index2 == 3189 || pixel_index2 == 3199 || pixel_index2 == 3245 || pixel_index2 == 3263 || pixel_index2 == 3266 || pixel_index2 == 3296 || pixel_index2 == 3332 || pixel_index2 == 3359 || pixel_index2 == 3362 || pixel_index2 == 3392 || pixel_index2 == 3440 || pixel_index2 == 3455 || pixel_index2 == 3458 || pixel_index2 == 3481 || pixel_index2 == 3488 || pixel_index2 == 3536 || pixel_index2 == 3551 || pixel_index2 == 3554 || ((pixel_index2 >= 3576) && (pixel_index2 <= 3577)) || pixel_index2 == 3583 || pixel_index2 == 3620 || pixel_index2 == 3632 || pixel_index2 == 3647 || pixel_index2 == 3650 || pixel_index2 == 3677 || pixel_index2 == 3718 || pixel_index2 == 3816 || ((pixel_index2 >= 3914) && (pixel_index2 <= 3918)) || pixel_index2 == 3937 || pixel_index2 == 4033 || pixel_index2 == 4129 || pixel_index2 == 4225 || pixel_index2 == 4317 || pixel_index2 == 4321 || pixel_index2 == 4413 || pixel_index2 == 4417 || pixel_index2 == 4703 || pixel_index2 == 4799 || pixel_index2 == 4895 || pixel_index2 == 4926 || pixel_index2 == 4930 || ((pixel_index2 >= 4956) && (pixel_index2 <= 4957)) || pixel_index2 == 4959 || pixel_index2 == 4991 || pixel_index2 == 5058 || pixel_index2 == 5087 || pixel_index2 == 5115 || pixel_index2 == 5211 || pixel_index2 == 5281 || pixel_index2 == 5307 || pixel_index2 == 5376 || pixel_index2 == 5403 || pixel_index2 == 5499 || pixel_index2 == 5585 || ((pixel_index2 >= 5587) && (pixel_index2 <= 5588)) || pixel_index2 == 5592 || pixel_index2 == 5679 || pixel_index2 == 5771 || pixel_index2 == 5810 || pixel_index2 == 5819 || ((pixel_index2 >= 5835) && (pixel_index2 <= 5836)) || pixel_index2 == 5866 || (pixel_index2 >= 5959) && (pixel_index2 <= 5962)) oled_data2 = 16'b0101001010000000;
        else if (pixel_index2 == 194 || pixel_index2 == 215 || pixel_index2 == 219 || pixel_index2 == 226 || pixel_index2 == 233 || pixel_index2 == 250 || pixel_index2 == 256 || pixel_index2 == 333 || pixel_index2 == 389 || pixel_index2 == 429 || ((pixel_index2 >= 509) && (pixel_index2 <= 510)) || pixel_index2 == 600 || pixel_index2 == 747 || pixel_index2 == 875 || pixel_index2 == 902 || pixel_index2 == 907 || pixel_index2 == 936 || ((pixel_index2 >= 968) && (pixel_index2 <= 969)) || pixel_index2 == 987 || pixel_index2 == 994 || pixel_index2 == 1001 || pixel_index2 == 1012 || pixel_index2 == 1019 || pixel_index2 == 1028 || pixel_index2 == 1031 || pixel_index2 == 1043 || ((pixel_index2 >= 5017) && (pixel_index2 <= 5018)) || ((pixel_index2 >= 5022) && (pixel_index2 <= 5023)) || pixel_index2 == 5026 || pixel_index2 == 5029 || pixel_index2 == 5036 || pixel_index2 == 5046 || pixel_index2 == 5049 || ((pixel_index2 >= 5052) && (pixel_index2 <= 5053)) || pixel_index2 == 5059 || pixel_index2 == 5063 || pixel_index2 == 5141 || pixel_index2 == 5245 || pixel_index2 == 5336 || pixel_index2 == 5629 || pixel_index2 == 5813) oled_data2 = 16'b1111011110010100;
        else if (pixel_index2 == 195 || ((pixel_index2 >= 200) && (pixel_index2 <= 201)) || ((pixel_index2 >= 206) && (pixel_index2 <= 207)) || ((pixel_index2 >= 210) && (pixel_index2 <= 212)) || pixel_index2 == 216 || pixel_index2 == 218 || pixel_index2 == 229 || pixel_index2 == 232 || ((pixel_index2 >= 238) && (pixel_index2 <= 240)) || ((pixel_index2 >= 243) && (pixel_index2 <= 244)) || pixel_index2 == 248 || pixel_index2 == 251 || pixel_index2 == 257 || ((pixel_index2 >= 259) && (pixel_index2 <= 260)) || ((pixel_index2 >= 263) && (pixel_index2 <= 264)) || pixel_index2 == 266 || ((pixel_index2 >= 269) && (pixel_index2 <= 272)) || pixel_index2 == 275 || ((pixel_index2 >= 278) && (pixel_index2 <= 279)) || ((pixel_index2 >= 284) && (pixel_index2 <= 285)) || ((pixel_index2 >= 290) && (pixel_index2 <= 291)) || ((pixel_index2 >= 296) && (pixel_index2 <= 297)) || ((pixel_index2 >= 302) && (pixel_index2 <= 303)) || ((pixel_index2 >= 306) && (pixel_index2 <= 308)) || ((pixel_index2 >= 311) && (pixel_index2 <= 312)) || ((pixel_index2 >= 314) && (pixel_index2 <= 315)) || pixel_index2 == 322 || ((pixel_index2 >= 325) && (pixel_index2 <= 326)) || ((pixel_index2 >= 328) && (pixel_index2 <= 329)) || ((pixel_index2 >= 334) && (pixel_index2 <= 336)) || ((pixel_index2 >= 338) && (pixel_index2 <= 340)) || ((pixel_index2 >= 343) && (pixel_index2 <= 344)) || pixel_index2 == 347 || ((pixel_index2 >= 352) && (pixel_index2 <= 353)) || ((pixel_index2 >= 355) && (pixel_index2 <= 356)) || pixel_index2 == 359 || ((pixel_index2 >= 362) && (pixel_index2 <= 363)) || ((pixel_index2 >= 367) && (pixel_index2 <= 368)) || pixel_index2 == 371 || ((pixel_index2 >= 374) && (pixel_index2 <= 375)) || ((pixel_index2 >= 380) && (pixel_index2 <= 381)) || ((pixel_index2 >= 386) && (pixel_index2 <= 387)) || pixel_index2 == 390 || ((pixel_index2 >= 392) && (pixel_index2 <= 393)) || ((pixel_index2 >= 397) && (pixel_index2 <= 400)) || ((pixel_index2 >= 402) && (pixel_index2 <= 404)) || ((pixel_index2 >= 407) && (pixel_index2 <= 408)) || pixel_index2 == 418 || ((pixel_index2 >= 421) && (pixel_index2 <= 422)) || ((pixel_index2 >= 424) && (pixel_index2 <= 425)) || pixel_index2 == 430 || pixel_index2 == 432 || pixel_index2 == 434 || pixel_index2 == 436 || ((pixel_index2 >= 439) && (pixel_index2 <= 440)) || ((pixel_index2 >= 448) && (pixel_index2 <= 449)) || pixel_index2 == 455 || ((pixel_index2 >= 463) && (pixel_index2 <= 464)) || pixel_index2 == 467 || ((pixel_index2 >= 470) && (pixel_index2 <= 471)) || ((pixel_index2 >= 476) && (pixel_index2 <= 477)) || ((pixel_index2 >= 482) && (pixel_index2 <= 483)) || ((pixel_index2 >= 488) && (pixel_index2 <= 489)) || ((pixel_index2 >= 493) && (pixel_index2 <= 494)) || pixel_index2 == 496 || pixel_index2 == 498 || pixel_index2 == 500 || ((pixel_index2 >= 503) && (pixel_index2 <= 504)) || pixel_index2 == 511 || pixel_index2 == 514 || ((pixel_index2 >= 517) && (pixel_index2 <= 518)) || ((pixel_index2 >= 520) && (pixel_index2 <= 521)) || ((pixel_index2 >= 525) && (pixel_index2 <= 526)) || pixel_index2 == 528 || pixel_index2 == 530 || ((pixel_index2 >= 532) && (pixel_index2 <= 533)) || ((pixel_index2 >= 536) && (pixel_index2 <= 537)) || ((pixel_index2 >= 544) && (pixel_index2 <= 546)) || ((pixel_index2 >= 551) && (pixel_index2 <= 552)) || ((pixel_index2 >= 559) && (pixel_index2 <= 560)) || pixel_index2 == 563 || ((pixel_index2 >= 566) && (pixel_index2 <= 567)) || ((pixel_index2 >= 572) && (pixel_index2 <= 573)) || ((pixel_index2 >= 578) && (pixel_index2 <= 579)) || pixel_index2 == 581 || ((pixel_index2 >= 584) && (pixel_index2 <= 585)) || ((pixel_index2 >= 589) && (pixel_index2 <= 590)) || pixel_index2 == 592 || pixel_index2 == 594 || pixel_index2 == 596 || ((pixel_index2 >= 601) && (pixel_index2 <= 602)) || pixel_index2 == 610 || ((pixel_index2 >= 613) && (pixel_index2 <= 614)) || ((pixel_index2 >= 616) && (pixel_index2 <= 617)) || ((pixel_index2 >= 621) && (pixel_index2 <= 622)) || pixel_index2 == 624 || pixel_index2 == 626 || ((pixel_index2 >= 628) && (pixel_index2 <= 629)) || ((pixel_index2 >= 633) && (pixel_index2 <= 634)) || ((pixel_index2 >= 641) && (pixel_index2 <= 643)) || ((pixel_index2 >= 648) && (pixel_index2 <= 650)) || ((pixel_index2 >= 653) && (pixel_index2 <= 656)) || ((pixel_index2 >= 660) && (pixel_index2 <= 663)) || ((pixel_index2 >= 666) && (pixel_index2 <= 669)) || ((pixel_index2 >= 674) && (pixel_index2 <= 675)) || pixel_index2 == 677 || ((pixel_index2 >= 680) && (pixel_index2 <= 681)) || ((pixel_index2 >= 685) && (pixel_index2 <= 686)) || ((pixel_index2 >= 688) && (pixel_index2 <= 690)) || pixel_index2 == 692 || ((pixel_index2 >= 698) && (pixel_index2 <= 699)) || pixel_index2 == 706 || ((pixel_index2 >= 709) && (pixel_index2 <= 710)) || ((pixel_index2 >= 712) && (pixel_index2 <= 713)) || ((pixel_index2 >= 717) && (pixel_index2 <= 718)) || ((pixel_index2 >= 720) && (pixel_index2 <= 722)) || ((pixel_index2 >= 724) && (pixel_index2 <= 725)) || ((pixel_index2 >= 730) && (pixel_index2 <= 731)) || ((pixel_index2 >= 739) && (pixel_index2 <= 740)) || pixel_index2 == 746 || ((pixel_index2 >= 751) && (pixel_index2 <= 752)) || pixel_index2 == 755 || ((pixel_index2 >= 758) && (pixel_index2 <= 759)) || ((pixel_index2 >= 761) && (pixel_index2 <= 762)) || ((pixel_index2 >= 764) && (pixel_index2 <= 765)) || ((pixel_index2 >= 770) && (pixel_index2 <= 771)) || ((pixel_index2 >= 776) && (pixel_index2 <= 777)) || ((pixel_index2 >= 781) && (pixel_index2 <= 782)) || ((pixel_index2 >= 784) && (pixel_index2 <= 786)) || ((pixel_index2 >= 788) && (pixel_index2 <= 789)) || ((pixel_index2 >= 794) && (pixel_index2 <= 795)) || pixel_index2 == 802 || ((pixel_index2 >= 805) && (pixel_index2 <= 806)) || ((pixel_index2 >= 808) && (pixel_index2 <= 809)) || ((pixel_index2 >= 813) && (pixel_index2 <= 814)) || ((pixel_index2 >= 816) && (pixel_index2 <= 818)) || ((pixel_index2 >= 820) && (pixel_index2 <= 821)) || pixel_index2 == 827 || ((pixel_index2 >= 835) && (pixel_index2 <= 836)) || ((pixel_index2 >= 842) && (pixel_index2 <= 843)) || ((pixel_index2 >= 847) && (pixel_index2 <= 848)) || pixel_index2 == 851 || ((pixel_index2 >= 854) && (pixel_index2 <= 855)) || ((pixel_index2 >= 857) && (pixel_index2 <= 858)) || ((pixel_index2 >= 860) && (pixel_index2 <= 861)) || ((pixel_index2 >= 866) && (pixel_index2 <= 868)) || ((pixel_index2 >= 872) && (pixel_index2 <= 874)) || ((pixel_index2 >= 877) && (pixel_index2 <= 878)) || ((pixel_index2 >= 880) && (pixel_index2 <= 881)) || ((pixel_index2 >= 884) && (pixel_index2 <= 885)) || ((pixel_index2 >= 887) && (pixel_index2 <= 888)) || ((pixel_index2 >= 890) && (pixel_index2 <= 891)) || pixel_index2 == 898 || pixel_index2 == 901 || ((pixel_index2 >= 904) && (pixel_index2 <= 906)) || ((pixel_index2 >= 909) && (pixel_index2 <= 910)) || ((pixel_index2 >= 912) && (pixel_index2 <= 914)) || ((pixel_index2 >= 916) && (pixel_index2 <= 917)) || pixel_index2 == 920 || pixel_index2 == 923 || ((pixel_index2 >= 928) && (pixel_index2 <= 929)) || ((pixel_index2 >= 931) && (pixel_index2 <= 932)) || pixel_index2 == 935 || ((pixel_index2 >= 938) && (pixel_index2 <= 939)) || ((pixel_index2 >= 943) && (pixel_index2 <= 944)) || pixel_index2 == 947 || ((pixel_index2 >= 950) && (pixel_index2 <= 951)) || ((pixel_index2 >= 953) && (pixel_index2 <= 954)) || ((pixel_index2 >= 956) && (pixel_index2 <= 957)) || ((pixel_index2 >= 962) && (pixel_index2 <= 964)) || pixel_index2 == 973 || ((pixel_index2 >= 976) && (pixel_index2 <= 977)) || ((pixel_index2 >= 980) && (pixel_index2 <= 981)) || ((pixel_index2 >= 984) && (pixel_index2 <= 986)) || ((pixel_index2 >= 995) && (pixel_index2 <= 997)) || pixel_index2 == 1000 || pixel_index2 == 1005 || ((pixel_index2 >= 1008) && (pixel_index2 <= 1010)) || pixel_index2 == 1013 || ((pixel_index2 >= 1016) && (pixel_index2 <= 1018)) || ((pixel_index2 >= 1025) && (pixel_index2 <= 1027)) || ((pixel_index2 >= 1032) && (pixel_index2 <= 1034)) || ((pixel_index2 >= 1037) && (pixel_index2 <= 1040)) || ((pixel_index2 >= 1044) && (pixel_index2 <= 1047)) || ((pixel_index2 >= 1050) && (pixel_index2 <= 1053)) || ((pixel_index2 >= 5030) && (pixel_index2 <= 5032)) || ((pixel_index2 >= 5037) && (pixel_index2 <= 5040)) || ((pixel_index2 >= 5047) && (pixel_index2 <= 5048)) || ((pixel_index2 >= 5055) && (pixel_index2 <= 5056)) || ((pixel_index2 >= 5060) && (pixel_index2 <= 5062)) || ((pixel_index2 >= 5113) && (pixel_index2 <= 5114)) || ((pixel_index2 >= 5118) && (pixel_index2 <= 5119)) || pixel_index2 == 5122 || ((pixel_index2 >= 5125) && (pixel_index2 <= 5126)) || ((pixel_index2 >= 5128) && (pixel_index2 <= 5129)) || ((pixel_index2 >= 5132) && (pixel_index2 <= 5133)) || ((pixel_index2 >= 5135) && (pixel_index2 <= 5136)) || pixel_index2 == 5142 || ((pixel_index2 >= 5144) && (pixel_index2 <= 5145)) || ((pixel_index2 >= 5148) && (pixel_index2 <= 5149)) || ((pixel_index2 >= 5151) && (pixel_index2 <= 5152)) || ((pixel_index2 >= 5155) && (pixel_index2 <= 5156)) || ((pixel_index2 >= 5158) && (pixel_index2 <= 5159)) || ((pixel_index2 >= 5209) && (pixel_index2 <= 5210)) || ((pixel_index2 >= 5214) && (pixel_index2 <= 5215)) || pixel_index2 == 5218 || ((pixel_index2 >= 5221) && (pixel_index2 <= 5222)) || ((pixel_index2 >= 5224) && (pixel_index2 <= 5225)) || pixel_index2 == 5228 || ((pixel_index2 >= 5231) && (pixel_index2 <= 5232)) || ((pixel_index2 >= 5237) && (pixel_index2 <= 5238)) || ((pixel_index2 >= 5240) && (pixel_index2 <= 5241)) || pixel_index2 == 5244 || ((pixel_index2 >= 5247) && (pixel_index2 <= 5248)) || ((pixel_index2 >= 5251) && (pixel_index2 <= 5252)) || ((pixel_index2 >= 5254) && (pixel_index2 <= 5255)) || ((pixel_index2 >= 5305) && (pixel_index2 <= 5306)) || ((pixel_index2 >= 5310) && (pixel_index2 <= 5312)) || pixel_index2 == 5314 || ((pixel_index2 >= 5317) && (pixel_index2 <= 5318)) || ((pixel_index2 >= 5320) && (pixel_index2 <= 5321)) || pixel_index2 == 5324 || ((pixel_index2 >= 5327) && (pixel_index2 <= 5328)) || ((pixel_index2 >= 5333) && (pixel_index2 <= 5334)) || pixel_index2 == 5337 || ((pixel_index2 >= 5340) && (pixel_index2 <= 5341)) || ((pixel_index2 >= 5343) && (pixel_index2 <= 5344)) || ((pixel_index2 >= 5347) && (pixel_index2 <= 5348)) || ((pixel_index2 >= 5350) && (pixel_index2 <= 5351)) || ((pixel_index2 >= 5401) && (pixel_index2 <= 5402)) || ((pixel_index2 >= 5406) && (pixel_index2 <= 5410)) || ((pixel_index2 >= 5413) && (pixel_index2 <= 5414)) || ((pixel_index2 >= 5416) && (pixel_index2 <= 5417)) || pixel_index2 == 5420 || ((pixel_index2 >= 5423) && (pixel_index2 <= 5424)) || ((pixel_index2 >= 5429) && (pixel_index2 <= 5430)) || ((pixel_index2 >= 5432) && (pixel_index2 <= 5433)) || pixel_index2 == 5437 || ((pixel_index2 >= 5439) && (pixel_index2 <= 5440)) || ((pixel_index2 >= 5443) && (pixel_index2 <= 5444)) || ((pixel_index2 >= 5446) && (pixel_index2 <= 5447)) || ((pixel_index2 >= 5497) && (pixel_index2 <= 5498)) || pixel_index2 == 5502 || ((pixel_index2 >= 5504) && (pixel_index2 <= 5506)) || ((pixel_index2 >= 5509) && (pixel_index2 <= 5510)) || ((pixel_index2 >= 5512) && (pixel_index2 <= 5513)) || pixel_index2 == 5516 || ((pixel_index2 >= 5519) && (pixel_index2 <= 5520)) || ((pixel_index2 >= 5525) && (pixel_index2 <= 5526)) || ((pixel_index2 >= 5528) && (pixel_index2 <= 5529)) || ((pixel_index2 >= 5533) && (pixel_index2 <= 5536)) || ((pixel_index2 >= 5540) && (pixel_index2 <= 5543)) || ((pixel_index2 >= 5593) && (pixel_index2 <= 5594)) || pixel_index2 == 5598 || ((pixel_index2 >= 5601) && (pixel_index2 <= 5602)) || ((pixel_index2 >= 5605) && (pixel_index2 <= 5606)) || ((pixel_index2 >= 5608) && (pixel_index2 <= 5609)) || pixel_index2 == 5612 || ((pixel_index2 >= 5615) && (pixel_index2 <= 5616)) || ((pixel_index2 >= 5621) && (pixel_index2 <= 5622)) || ((pixel_index2 >= 5624) && (pixel_index2 <= 5625)) || pixel_index2 == 5628 || ((pixel_index2 >= 5631) && (pixel_index2 <= 5632)) || ((pixel_index2 >= 5635) && (pixel_index2 <= 5636)) || ((pixel_index2 >= 5638) && (pixel_index2 <= 5639)) || ((pixel_index2 >= 5689) && (pixel_index2 <= 5690)) || pixel_index2 == 5694 || ((pixel_index2 >= 5697) && (pixel_index2 <= 5698)) || ((pixel_index2 >= 5701) && (pixel_index2 <= 5702)) || ((pixel_index2 >= 5704) && (pixel_index2 <= 5705)) || pixel_index2 == 5708 || ((pixel_index2 >= 5711) && (pixel_index2 <= 5712)) || ((pixel_index2 >= 5717) && (pixel_index2 <= 5718)) || ((pixel_index2 >= 5720) && (pixel_index2 <= 5721)) || ((pixel_index2 >= 5724) && (pixel_index2 <= 5725)) || ((pixel_index2 >= 5727) && (pixel_index2 <= 5728)) || ((pixel_index2 >= 5731) && (pixel_index2 <= 5732)) || ((pixel_index2 >= 5734) && (pixel_index2 <= 5735)) || ((pixel_index2 >= 5783) && (pixel_index2 <= 5787)) || pixel_index2 == 5790 || ((pixel_index2 >= 5793) && (pixel_index2 <= 5794)) || ((pixel_index2 >= 5797) && (pixel_index2 <= 5798)) || ((pixel_index2 >= 5800) && (pixel_index2 <= 5801)) || ((pixel_index2 >= 5804) && (pixel_index2 <= 5805)) || ((pixel_index2 >= 5807) && (pixel_index2 <= 5808)) || pixel_index2 == 5814 || ((pixel_index2 >= 5816) && (pixel_index2 <= 5817)) || ((pixel_index2 >= 5820) && (pixel_index2 <= 5821)) || ((pixel_index2 >= 5823) && (pixel_index2 <= 5824)) || ((pixel_index2 >= 5827) && (pixel_index2 <= 5828)) || ((pixel_index2 >= 5830) && (pixel_index2 <= 5831)) || pixel_index2 == 5895 || pixel_index2 == 5911) oled_data2 = 16'b1111011110011110;
        else if (pixel_index2 == 227 || pixel_index2 == 301 || pixel_index2 == 435 || pixel_index2 == 437 || pixel_index2 == 485 || pixel_index2 == 505 || pixel_index2 == 593 || pixel_index2 == 665 || pixel_index2 == 745 || pixel_index2 == 5912) oled_data2 = 16'b1010011110010100;
        else if (pixel_index2 == 900) oled_data2 = 16'b0101010100001010;
        else if (pixel_index2 == 5972 || pixel_index2 == 5974 || pixel_index2 == 6062 || pixel_index2 == 6064 || (pixel_index2 >= 6068) && (pixel_index2 <= 6070)) oled_data2 = 16'b0000000000001010;
        else if (pixel_index2 == 6059) oled_data2 = 16'b0000001010000000;
        else if (pixel_index2 == 6063) oled_data2 = 16'b0000001010001010;
        else oled_data2 = 0;
    end
end

endmodule 