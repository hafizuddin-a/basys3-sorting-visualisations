`timescale 1ns / 1ps

module selection_sort(

    );
endmodule
